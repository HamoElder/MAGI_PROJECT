// Generator : SpinalHDL v1.7.0    git head : eca519e78d4e6022e34911ec300a432ed9db8220
// Component : AxiLite4MIMOReceiver
// Git hash  : a61652a25e7e73fd6a89f26f1edce017e805a730

`timescale 1ns/1ps

module AxiLite4MIMOReceiver (
  input               axil4Ctrl_awvalid,
  output              axil4Ctrl_awready,
  input      [7:0]    axil4Ctrl_awaddr,
  input      [2:0]    axil4Ctrl_awprot,
  input               axil4Ctrl_wvalid,
  output              axil4Ctrl_wready,
  input      [31:0]   axil4Ctrl_wdata,
  input      [3:0]    axil4Ctrl_wstrb,
  output              axil4Ctrl_bvalid,
  input               axil4Ctrl_bready,
  output     [1:0]    axil4Ctrl_bresp,
  input               axil4Ctrl_arvalid,
  output reg          axil4Ctrl_arready,
  input      [7:0]    axil4Ctrl_araddr,
  input      [2:0]    axil4Ctrl_arprot,
  output              axil4Ctrl_rvalid,
  input               axil4Ctrl_rready,
  output     [31:0]   axil4Ctrl_rdata,
  output     [1:0]    axil4Ctrl_rresp,
  input               mod_iq_valid,
  output              mod_iq_ready,
  input      [15:0]   mod_iq_payload_cha_i,
  input      [15:0]   mod_iq_payload_cha_q,
  output              base_sub_iqs_valid,
  output     [31:0]   base_sub_iqs_payload_0_cha_i,
  output     [31:0]   base_sub_iqs_payload_0_cha_q,
  output     [31:0]   base_sub_iqs_payload_1_cha_i,
  output     [31:0]   base_sub_iqs_payload_1_cha_q,
  output     [31:0]   base_sub_iqs_payload_2_cha_i,
  output     [31:0]   base_sub_iqs_payload_2_cha_q,
  output     [31:0]   base_sub_iqs_payload_3_cha_i,
  output     [31:0]   base_sub_iqs_payload_3_cha_q,
  output     [31:0]   base_sub_iqs_payload_4_cha_i,
  output     [31:0]   base_sub_iqs_payload_4_cha_q,
  output     [31:0]   base_sub_iqs_payload_5_cha_i,
  output     [31:0]   base_sub_iqs_payload_5_cha_q,
  output     [31:0]   base_sub_iqs_payload_6_cha_i,
  output     [31:0]   base_sub_iqs_payload_6_cha_q,
  output     [31:0]   base_sub_iqs_payload_7_cha_i,
  output     [31:0]   base_sub_iqs_payload_7_cha_q,
  input               rf_clk,
  input               rf_resetn,
  input               clk,
  input               resetn
);

  wire                rfClockArea_mimo_receiver_mod_iq_ready;
  wire                rfClockArea_mimo_receiver_base_sub_iqs_valid;
  wire       [31:0]   rfClockArea_mimo_receiver_base_sub_iqs_payload_0_cha_i;
  wire       [31:0]   rfClockArea_mimo_receiver_base_sub_iqs_payload_0_cha_q;
  wire       [31:0]   rfClockArea_mimo_receiver_base_sub_iqs_payload_1_cha_i;
  wire       [31:0]   rfClockArea_mimo_receiver_base_sub_iqs_payload_1_cha_q;
  wire       [31:0]   rfClockArea_mimo_receiver_base_sub_iqs_payload_2_cha_i;
  wire       [31:0]   rfClockArea_mimo_receiver_base_sub_iqs_payload_2_cha_q;
  wire       [31:0]   rfClockArea_mimo_receiver_base_sub_iqs_payload_3_cha_i;
  wire       [31:0]   rfClockArea_mimo_receiver_base_sub_iqs_payload_3_cha_q;
  wire       [31:0]   rfClockArea_mimo_receiver_base_sub_iqs_payload_4_cha_i;
  wire       [31:0]   rfClockArea_mimo_receiver_base_sub_iqs_payload_4_cha_q;
  wire       [31:0]   rfClockArea_mimo_receiver_base_sub_iqs_payload_5_cha_i;
  wire       [31:0]   rfClockArea_mimo_receiver_base_sub_iqs_payload_5_cha_q;
  wire       [31:0]   rfClockArea_mimo_receiver_base_sub_iqs_payload_6_cha_i;
  wire       [31:0]   rfClockArea_mimo_receiver_base_sub_iqs_payload_6_cha_q;
  wire       [31:0]   rfClockArea_mimo_receiver_base_sub_iqs_payload_7_cha_i;
  wire       [31:0]   rfClockArea_mimo_receiver_base_sub_iqs_payload_7_cha_q;
  wire                clkCrossing_4_dataOut;
  wire                clkCrossing_5_dataOut;
  wire       [5:0]    clkCrossing_6_dataOut;
  wire       [15:0]   clkCrossing_7_dataOut;
  wire                readHaltRequest;
  wire                writeHaltRequest;
  wire                writeJoinEvent_valid;
  wire                writeJoinEvent_ready;
  wire                writeJoinEvent_fire;
  wire       [1:0]    writeRsp_resp;
  wire                writeJoinEvent_translated_valid;
  wire                writeJoinEvent_translated_ready;
  wire       [1:0]    writeJoinEvent_translated_payload_resp;
  wire                _zz_axil4Ctrl_bvalid;
  reg                 _zz_writeJoinEvent_translated_ready;
  wire                _zz_axil4Ctrl_bvalid_1;
  reg                 _zz_axil4Ctrl_bvalid_2;
  reg        [1:0]    _zz_axil4Ctrl_bresp;
  wire                when_Stream_l368;
  wire                readDataStage_valid;
  wire                readDataStage_ready;
  wire       [7:0]    readDataStage_payload_addr;
  wire       [2:0]    readDataStage_payload_prot;
  reg                 axil4Ctrl_ar_rValid;
  reg        [7:0]    axil4Ctrl_ar_rData_addr;
  reg        [2:0]    axil4Ctrl_ar_rData_prot;
  wire                when_Stream_l368_1;
  reg        [31:0]   readRsp_data;
  wire       [1:0]    readRsp_resp;
  wire                _zz_axil4Ctrl_rvalid;
  wire                writeOccur;
  wire                readOccur;
  wire                oam_unspinor_bridge_w_sel;
  wire                oam_unspinor_bridge_w_en;
  wire       [5:0]    oam_unspinor_bridge_w_addr;
  wire       [15:0]   oam_unspinor_bridge_w_data;
  reg                 oam_unspinor_bridge_w_en_driver;
  reg                 oam_unspinor_bridge_w_sel_driver;
  reg        [5:0]    _zz_oam_unspinor_bridge_w_addr;
  reg        [15:0]   _zz_oam_unspinor_bridge_w_data;

  MIMOReceiver rfClockArea_mimo_receiver (
    .mod_iq_valid                 (mod_iq_valid                                                ), //i
    .mod_iq_ready                 (rfClockArea_mimo_receiver_mod_iq_ready                      ), //o
    .mod_iq_payload_cha_i         (mod_iq_payload_cha_i[15:0]                                  ), //i
    .mod_iq_payload_cha_q         (mod_iq_payload_cha_q[15:0]                                  ), //i
    .base_sub_iqs_valid           (rfClockArea_mimo_receiver_base_sub_iqs_valid                ), //o
    .base_sub_iqs_payload_0_cha_i (rfClockArea_mimo_receiver_base_sub_iqs_payload_0_cha_i[31:0]), //o
    .base_sub_iqs_payload_0_cha_q (rfClockArea_mimo_receiver_base_sub_iqs_payload_0_cha_q[31:0]), //o
    .base_sub_iqs_payload_1_cha_i (rfClockArea_mimo_receiver_base_sub_iqs_payload_1_cha_i[31:0]), //o
    .base_sub_iqs_payload_1_cha_q (rfClockArea_mimo_receiver_base_sub_iqs_payload_1_cha_q[31:0]), //o
    .base_sub_iqs_payload_2_cha_i (rfClockArea_mimo_receiver_base_sub_iqs_payload_2_cha_i[31:0]), //o
    .base_sub_iqs_payload_2_cha_q (rfClockArea_mimo_receiver_base_sub_iqs_payload_2_cha_q[31:0]), //o
    .base_sub_iqs_payload_3_cha_i (rfClockArea_mimo_receiver_base_sub_iqs_payload_3_cha_i[31:0]), //o
    .base_sub_iqs_payload_3_cha_q (rfClockArea_mimo_receiver_base_sub_iqs_payload_3_cha_q[31:0]), //o
    .base_sub_iqs_payload_4_cha_i (rfClockArea_mimo_receiver_base_sub_iqs_payload_4_cha_i[31:0]), //o
    .base_sub_iqs_payload_4_cha_q (rfClockArea_mimo_receiver_base_sub_iqs_payload_4_cha_q[31:0]), //o
    .base_sub_iqs_payload_5_cha_i (rfClockArea_mimo_receiver_base_sub_iqs_payload_5_cha_i[31:0]), //o
    .base_sub_iqs_payload_5_cha_q (rfClockArea_mimo_receiver_base_sub_iqs_payload_5_cha_q[31:0]), //o
    .base_sub_iqs_payload_6_cha_i (rfClockArea_mimo_receiver_base_sub_iqs_payload_6_cha_i[31:0]), //o
    .base_sub_iqs_payload_6_cha_q (rfClockArea_mimo_receiver_base_sub_iqs_payload_6_cha_q[31:0]), //o
    .base_sub_iqs_payload_7_cha_i (rfClockArea_mimo_receiver_base_sub_iqs_payload_7_cha_i[31:0]), //o
    .base_sub_iqs_payload_7_cha_q (rfClockArea_mimo_receiver_base_sub_iqs_payload_7_cha_q[31:0]), //o
    .w_sel                        (clkCrossing_5_dataOut                                       ), //i
    .w_en                         (clkCrossing_4_dataOut                                       ), //i
    .w_addr                       (clkCrossing_6_dataOut[5:0]                                  ), //i
    .w_data                       (clkCrossing_7_dataOut[15:0]                                 ), //i
    .rf_clk                       (rf_clk                                                      ), //i
    .rf_resetn                    (rf_resetn                                                   )  //i
  );
  ClkCrossing clkCrossing_4 (
    .dataIn    (oam_unspinor_bridge_w_en), //i
    .dataOut   (clkCrossing_4_dataOut   ), //o
    .clk       (clk                     ), //i
    .resetn    (resetn                  ), //i
    .rf_clk    (rf_clk                  ), //i
    .rf_resetn (rf_resetn               )  //i
  );
  ClkCrossing clkCrossing_5 (
    .dataIn    (oam_unspinor_bridge_w_sel), //i
    .dataOut   (clkCrossing_5_dataOut    ), //o
    .clk       (clk                      ), //i
    .resetn    (resetn                   ), //i
    .rf_clk    (rf_clk                   ), //i
    .rf_resetn (rf_resetn                )  //i
  );
  ClkCrossing_2 clkCrossing_6 (
    .dataIn    (oam_unspinor_bridge_w_addr[5:0]), //i
    .dataOut   (clkCrossing_6_dataOut[5:0]     ), //o
    .clk       (clk                            ), //i
    .resetn    (resetn                         ), //i
    .rf_clk    (rf_clk                         ), //i
    .rf_resetn (rf_resetn                      )  //i
  );
  ClkCrossing_3 clkCrossing_7 (
    .dataIn    (oam_unspinor_bridge_w_data[15:0]), //i
    .dataOut   (clkCrossing_7_dataOut[15:0]     ), //o
    .clk       (clk                             ), //i
    .resetn    (resetn                          ), //i
    .rf_clk    (rf_clk                          ), //i
    .rf_resetn (rf_resetn                       )  //i
  );
  assign mod_iq_ready = rfClockArea_mimo_receiver_mod_iq_ready;
  assign base_sub_iqs_valid = rfClockArea_mimo_receiver_base_sub_iqs_valid;
  assign base_sub_iqs_payload_0_cha_i = rfClockArea_mimo_receiver_base_sub_iqs_payload_0_cha_i;
  assign base_sub_iqs_payload_0_cha_q = rfClockArea_mimo_receiver_base_sub_iqs_payload_0_cha_q;
  assign base_sub_iqs_payload_1_cha_i = rfClockArea_mimo_receiver_base_sub_iqs_payload_1_cha_i;
  assign base_sub_iqs_payload_1_cha_q = rfClockArea_mimo_receiver_base_sub_iqs_payload_1_cha_q;
  assign base_sub_iqs_payload_2_cha_i = rfClockArea_mimo_receiver_base_sub_iqs_payload_2_cha_i;
  assign base_sub_iqs_payload_2_cha_q = rfClockArea_mimo_receiver_base_sub_iqs_payload_2_cha_q;
  assign base_sub_iqs_payload_3_cha_i = rfClockArea_mimo_receiver_base_sub_iqs_payload_3_cha_i;
  assign base_sub_iqs_payload_3_cha_q = rfClockArea_mimo_receiver_base_sub_iqs_payload_3_cha_q;
  assign base_sub_iqs_payload_4_cha_i = rfClockArea_mimo_receiver_base_sub_iqs_payload_4_cha_i;
  assign base_sub_iqs_payload_4_cha_q = rfClockArea_mimo_receiver_base_sub_iqs_payload_4_cha_q;
  assign base_sub_iqs_payload_5_cha_i = rfClockArea_mimo_receiver_base_sub_iqs_payload_5_cha_i;
  assign base_sub_iqs_payload_5_cha_q = rfClockArea_mimo_receiver_base_sub_iqs_payload_5_cha_q;
  assign base_sub_iqs_payload_6_cha_i = rfClockArea_mimo_receiver_base_sub_iqs_payload_6_cha_i;
  assign base_sub_iqs_payload_6_cha_q = rfClockArea_mimo_receiver_base_sub_iqs_payload_6_cha_q;
  assign base_sub_iqs_payload_7_cha_i = rfClockArea_mimo_receiver_base_sub_iqs_payload_7_cha_i;
  assign base_sub_iqs_payload_7_cha_q = rfClockArea_mimo_receiver_base_sub_iqs_payload_7_cha_q;
  assign readHaltRequest = 1'b0;
  assign writeHaltRequest = 1'b0;
  assign writeJoinEvent_fire = (writeJoinEvent_valid && writeJoinEvent_ready);
  assign writeJoinEvent_valid = (axil4Ctrl_awvalid && axil4Ctrl_wvalid);
  assign axil4Ctrl_awready = writeJoinEvent_fire;
  assign axil4Ctrl_wready = writeJoinEvent_fire;
  assign writeJoinEvent_translated_valid = writeJoinEvent_valid;
  assign writeJoinEvent_ready = writeJoinEvent_translated_ready;
  assign writeJoinEvent_translated_payload_resp = writeRsp_resp;
  assign _zz_axil4Ctrl_bvalid = (! writeHaltRequest);
  assign writeJoinEvent_translated_ready = (_zz_writeJoinEvent_translated_ready && _zz_axil4Ctrl_bvalid);
  always @(*) begin
    _zz_writeJoinEvent_translated_ready = axil4Ctrl_bready;
    if(when_Stream_l368) begin
      _zz_writeJoinEvent_translated_ready = 1'b1;
    end
  end

  assign when_Stream_l368 = (! _zz_axil4Ctrl_bvalid_1);
  assign _zz_axil4Ctrl_bvalid_1 = _zz_axil4Ctrl_bvalid_2;
  assign axil4Ctrl_bvalid = _zz_axil4Ctrl_bvalid_1;
  assign axil4Ctrl_bresp = _zz_axil4Ctrl_bresp;
  always @(*) begin
    axil4Ctrl_arready = readDataStage_ready;
    if(when_Stream_l368_1) begin
      axil4Ctrl_arready = 1'b1;
    end
  end

  assign when_Stream_l368_1 = (! readDataStage_valid);
  assign readDataStage_valid = axil4Ctrl_ar_rValid;
  assign readDataStage_payload_addr = axil4Ctrl_ar_rData_addr;
  assign readDataStage_payload_prot = axil4Ctrl_ar_rData_prot;
  assign _zz_axil4Ctrl_rvalid = (! readHaltRequest);
  assign readDataStage_ready = (axil4Ctrl_rready && _zz_axil4Ctrl_rvalid);
  assign axil4Ctrl_rvalid = (readDataStage_valid && _zz_axil4Ctrl_rvalid);
  assign axil4Ctrl_rdata = readRsp_data;
  assign axil4Ctrl_rresp = readRsp_resp;
  assign writeRsp_resp = 2'b00;
  assign readRsp_resp = 2'b00;
  always @(*) begin
    readRsp_data = 32'h0;
    case(readDataStage_payload_addr)
      8'h0 : begin
        readRsp_data[0 : 0] = oam_unspinor_bridge_w_en_driver;
        readRsp_data[1 : 1] = oam_unspinor_bridge_w_sel_driver;
      end
      default : begin
      end
    endcase
  end

  assign writeOccur = (writeJoinEvent_valid && writeJoinEvent_ready);
  assign readOccur = (axil4Ctrl_rvalid && axil4Ctrl_rready);
  assign oam_unspinor_bridge_w_en = oam_unspinor_bridge_w_en_driver;
  assign oam_unspinor_bridge_w_sel = oam_unspinor_bridge_w_sel_driver;
  assign oam_unspinor_bridge_w_addr = _zz_oam_unspinor_bridge_w_addr;
  assign oam_unspinor_bridge_w_data = _zz_oam_unspinor_bridge_w_data;
  always @(posedge clk) begin
    if(!resetn) begin
      _zz_axil4Ctrl_bvalid_2 <= 1'b0;
      axil4Ctrl_ar_rValid <= 1'b0;
      oam_unspinor_bridge_w_en_driver <= 1'b0;
      oam_unspinor_bridge_w_sel_driver <= 1'b0;
    end else begin
      if(_zz_writeJoinEvent_translated_ready) begin
        _zz_axil4Ctrl_bvalid_2 <= (writeJoinEvent_translated_valid && _zz_axil4Ctrl_bvalid);
      end
      if(axil4Ctrl_arready) begin
        axil4Ctrl_ar_rValid <= axil4Ctrl_arvalid;
      end
      case(axil4Ctrl_awaddr)
        8'h0 : begin
          if(writeOccur) begin
            oam_unspinor_bridge_w_en_driver <= axil4Ctrl_wdata[0];
            oam_unspinor_bridge_w_sel_driver <= axil4Ctrl_wdata[1];
          end
        end
        default : begin
        end
      endcase
    end
  end

  always @(posedge clk) begin
    if(_zz_writeJoinEvent_translated_ready) begin
      _zz_axil4Ctrl_bresp <= writeJoinEvent_translated_payload_resp;
    end
    if(axil4Ctrl_arready) begin
      axil4Ctrl_ar_rData_addr <= axil4Ctrl_araddr;
      axil4Ctrl_ar_rData_prot <= axil4Ctrl_arprot;
    end
    case(axil4Ctrl_awaddr)
      8'h04 : begin
        if(writeOccur) begin
          _zz_oam_unspinor_bridge_w_addr <= axil4Ctrl_wdata[5 : 0];
        end
      end
      8'h08 : begin
        if(writeOccur) begin
          _zz_oam_unspinor_bridge_w_data <= axil4Ctrl_wdata[15 : 0];
        end
      end
      default : begin
      end
    endcase
  end


endmodule

module ClkCrossing_3 (
  input      [15:0]   dataIn,
  output     [15:0]   dataOut,
  input               clk,
  input               resetn,
  input               rf_clk,
  input               rf_resetn
);

  reg        [15:0]   area_clkI_reg;
  (* async_reg = "true" *) reg        [15:0]   area_clkO_buf0;
  reg        [15:0]   area_clkO_buf1;

  assign dataOut = area_clkO_buf1;
  always @(posedge clk) begin
    area_clkI_reg <= dataIn;
  end

  always @(posedge rf_clk) begin
    area_clkO_buf0 <= area_clkI_reg;
    area_clkO_buf1 <= area_clkO_buf0;
  end


endmodule

module ClkCrossing_2 (
  input      [5:0]    dataIn,
  output     [5:0]    dataOut,
  input               clk,
  input               resetn,
  input               rf_clk,
  input               rf_resetn
);

  reg        [5:0]    area_clkI_reg;
  (* async_reg = "true" *) reg        [5:0]    area_clkO_buf0;
  reg        [5:0]    area_clkO_buf1;

  assign dataOut = area_clkO_buf1;
  always @(posedge clk) begin
    area_clkI_reg <= dataIn;
  end

  always @(posedge rf_clk) begin
    area_clkO_buf0 <= area_clkI_reg;
    area_clkO_buf1 <= area_clkO_buf0;
  end


endmodule

//ClkCrossing replaced by ClkCrossing

module ClkCrossing (
  input               dataIn,
  output              dataOut,
  input               clk,
  input               resetn,
  input               rf_clk,
  input               rf_resetn
);

  reg                 area_clkI_reg;
  (* async_reg = "true" *) reg                 area_clkO_buf0;
  reg                 area_clkO_buf1;

  assign dataOut = area_clkO_buf1;
  always @(posedge clk) begin
    area_clkI_reg <= dataIn;
  end

  always @(posedge rf_clk) begin
    area_clkO_buf0 <= area_clkI_reg;
    area_clkO_buf1 <= area_clkO_buf0;
  end


endmodule

module MIMOReceiver (
  input               mod_iq_valid,
  output              mod_iq_ready,
  input      [15:0]   mod_iq_payload_cha_i,
  input      [15:0]   mod_iq_payload_cha_q,
  output              base_sub_iqs_valid,
  output     [31:0]   base_sub_iqs_payload_0_cha_i,
  output     [31:0]   base_sub_iqs_payload_0_cha_q,
  output     [31:0]   base_sub_iqs_payload_1_cha_i,
  output     [31:0]   base_sub_iqs_payload_1_cha_q,
  output     [31:0]   base_sub_iqs_payload_2_cha_i,
  output     [31:0]   base_sub_iqs_payload_2_cha_q,
  output     [31:0]   base_sub_iqs_payload_3_cha_i,
  output     [31:0]   base_sub_iqs_payload_3_cha_q,
  output     [31:0]   base_sub_iqs_payload_4_cha_i,
  output     [31:0]   base_sub_iqs_payload_4_cha_q,
  output     [31:0]   base_sub_iqs_payload_5_cha_i,
  output     [31:0]   base_sub_iqs_payload_5_cha_q,
  output     [31:0]   base_sub_iqs_payload_6_cha_i,
  output     [31:0]   base_sub_iqs_payload_6_cha_q,
  output     [31:0]   base_sub_iqs_payload_7_cha_i,
  output     [31:0]   base_sub_iqs_payload_7_cha_q,
  input               w_sel,
  input               w_en,
  input      [5:0]    w_addr,
  input      [15:0]   w_data,
  input               rf_clk,
  input               rf_resetn
);

  wire       [15:0]   mIMOReceiverUnit_8_shift_i_0;
  wire       [15:0]   mIMOReceiverUnit_8_shift_i_1;
  wire       [15:0]   mIMOReceiverUnit_8_shift_i_2;
  wire       [15:0]   mIMOReceiverUnit_8_shift_i_3;
  wire       [15:0]   mIMOReceiverUnit_8_shift_i_4;
  wire       [15:0]   mIMOReceiverUnit_8_shift_i_5;
  wire       [15:0]   mIMOReceiverUnit_8_shift_i_6;
  wire       [15:0]   mIMOReceiverUnit_8_shift_i_7;
  wire       [15:0]   mIMOReceiverUnit_8_shift_q_0;
  wire       [15:0]   mIMOReceiverUnit_8_shift_q_1;
  wire       [15:0]   mIMOReceiverUnit_8_shift_q_2;
  wire       [15:0]   mIMOReceiverUnit_8_shift_q_3;
  wire       [15:0]   mIMOReceiverUnit_8_shift_q_4;
  wire       [15:0]   mIMOReceiverUnit_8_shift_q_5;
  wire       [15:0]   mIMOReceiverUnit_8_shift_q_6;
  wire       [15:0]   mIMOReceiverUnit_8_shift_q_7;
  wire       [15:0]   mIMOReceiverUnit_9_shift_i_0;
  wire       [15:0]   mIMOReceiverUnit_9_shift_i_1;
  wire       [15:0]   mIMOReceiverUnit_9_shift_i_2;
  wire       [15:0]   mIMOReceiverUnit_9_shift_i_3;
  wire       [15:0]   mIMOReceiverUnit_9_shift_i_4;
  wire       [15:0]   mIMOReceiverUnit_9_shift_i_5;
  wire       [15:0]   mIMOReceiverUnit_9_shift_i_6;
  wire       [15:0]   mIMOReceiverUnit_9_shift_i_7;
  wire       [15:0]   mIMOReceiverUnit_9_shift_q_0;
  wire       [15:0]   mIMOReceiverUnit_9_shift_q_1;
  wire       [15:0]   mIMOReceiverUnit_9_shift_q_2;
  wire       [15:0]   mIMOReceiverUnit_9_shift_q_3;
  wire       [15:0]   mIMOReceiverUnit_9_shift_q_4;
  wire       [15:0]   mIMOReceiverUnit_9_shift_q_5;
  wire       [15:0]   mIMOReceiverUnit_9_shift_q_6;
  wire       [15:0]   mIMOReceiverUnit_9_shift_q_7;
  wire       [15:0]   mIMOReceiverUnit_10_shift_i_0;
  wire       [15:0]   mIMOReceiverUnit_10_shift_i_1;
  wire       [15:0]   mIMOReceiverUnit_10_shift_i_2;
  wire       [15:0]   mIMOReceiverUnit_10_shift_i_3;
  wire       [15:0]   mIMOReceiverUnit_10_shift_i_4;
  wire       [15:0]   mIMOReceiverUnit_10_shift_i_5;
  wire       [15:0]   mIMOReceiverUnit_10_shift_i_6;
  wire       [15:0]   mIMOReceiverUnit_10_shift_i_7;
  wire       [15:0]   mIMOReceiverUnit_10_shift_q_0;
  wire       [15:0]   mIMOReceiverUnit_10_shift_q_1;
  wire       [15:0]   mIMOReceiverUnit_10_shift_q_2;
  wire       [15:0]   mIMOReceiverUnit_10_shift_q_3;
  wire       [15:0]   mIMOReceiverUnit_10_shift_q_4;
  wire       [15:0]   mIMOReceiverUnit_10_shift_q_5;
  wire       [15:0]   mIMOReceiverUnit_10_shift_q_6;
  wire       [15:0]   mIMOReceiverUnit_10_shift_q_7;
  wire       [15:0]   mIMOReceiverUnit_11_shift_i_0;
  wire       [15:0]   mIMOReceiverUnit_11_shift_i_1;
  wire       [15:0]   mIMOReceiverUnit_11_shift_i_2;
  wire       [15:0]   mIMOReceiverUnit_11_shift_i_3;
  wire       [15:0]   mIMOReceiverUnit_11_shift_i_4;
  wire       [15:0]   mIMOReceiverUnit_11_shift_i_5;
  wire       [15:0]   mIMOReceiverUnit_11_shift_i_6;
  wire       [15:0]   mIMOReceiverUnit_11_shift_i_7;
  wire       [15:0]   mIMOReceiverUnit_11_shift_q_0;
  wire       [15:0]   mIMOReceiverUnit_11_shift_q_1;
  wire       [15:0]   mIMOReceiverUnit_11_shift_q_2;
  wire       [15:0]   mIMOReceiverUnit_11_shift_q_3;
  wire       [15:0]   mIMOReceiverUnit_11_shift_q_4;
  wire       [15:0]   mIMOReceiverUnit_11_shift_q_5;
  wire       [15:0]   mIMOReceiverUnit_11_shift_q_6;
  wire       [15:0]   mIMOReceiverUnit_11_shift_q_7;
  wire       [15:0]   mIMOReceiverUnit_12_shift_i_0;
  wire       [15:0]   mIMOReceiverUnit_12_shift_i_1;
  wire       [15:0]   mIMOReceiverUnit_12_shift_i_2;
  wire       [15:0]   mIMOReceiverUnit_12_shift_i_3;
  wire       [15:0]   mIMOReceiverUnit_12_shift_i_4;
  wire       [15:0]   mIMOReceiverUnit_12_shift_i_5;
  wire       [15:0]   mIMOReceiverUnit_12_shift_i_6;
  wire       [15:0]   mIMOReceiverUnit_12_shift_i_7;
  wire       [15:0]   mIMOReceiverUnit_12_shift_q_0;
  wire       [15:0]   mIMOReceiverUnit_12_shift_q_1;
  wire       [15:0]   mIMOReceiverUnit_12_shift_q_2;
  wire       [15:0]   mIMOReceiverUnit_12_shift_q_3;
  wire       [15:0]   mIMOReceiverUnit_12_shift_q_4;
  wire       [15:0]   mIMOReceiverUnit_12_shift_q_5;
  wire       [15:0]   mIMOReceiverUnit_12_shift_q_6;
  wire       [15:0]   mIMOReceiverUnit_12_shift_q_7;
  wire       [15:0]   mIMOReceiverUnit_13_shift_i_0;
  wire       [15:0]   mIMOReceiverUnit_13_shift_i_1;
  wire       [15:0]   mIMOReceiverUnit_13_shift_i_2;
  wire       [15:0]   mIMOReceiverUnit_13_shift_i_3;
  wire       [15:0]   mIMOReceiverUnit_13_shift_i_4;
  wire       [15:0]   mIMOReceiverUnit_13_shift_i_5;
  wire       [15:0]   mIMOReceiverUnit_13_shift_i_6;
  wire       [15:0]   mIMOReceiverUnit_13_shift_i_7;
  wire       [15:0]   mIMOReceiverUnit_13_shift_q_0;
  wire       [15:0]   mIMOReceiverUnit_13_shift_q_1;
  wire       [15:0]   mIMOReceiverUnit_13_shift_q_2;
  wire       [15:0]   mIMOReceiverUnit_13_shift_q_3;
  wire       [15:0]   mIMOReceiverUnit_13_shift_q_4;
  wire       [15:0]   mIMOReceiverUnit_13_shift_q_5;
  wire       [15:0]   mIMOReceiverUnit_13_shift_q_6;
  wire       [15:0]   mIMOReceiverUnit_13_shift_q_7;
  wire       [15:0]   mIMOReceiverUnit_14_shift_i_0;
  wire       [15:0]   mIMOReceiverUnit_14_shift_i_1;
  wire       [15:0]   mIMOReceiverUnit_14_shift_i_2;
  wire       [15:0]   mIMOReceiverUnit_14_shift_i_3;
  wire       [15:0]   mIMOReceiverUnit_14_shift_i_4;
  wire       [15:0]   mIMOReceiverUnit_14_shift_i_5;
  wire       [15:0]   mIMOReceiverUnit_14_shift_i_6;
  wire       [15:0]   mIMOReceiverUnit_14_shift_i_7;
  wire       [15:0]   mIMOReceiverUnit_14_shift_q_0;
  wire       [15:0]   mIMOReceiverUnit_14_shift_q_1;
  wire       [15:0]   mIMOReceiverUnit_14_shift_q_2;
  wire       [15:0]   mIMOReceiverUnit_14_shift_q_3;
  wire       [15:0]   mIMOReceiverUnit_14_shift_q_4;
  wire       [15:0]   mIMOReceiverUnit_14_shift_q_5;
  wire       [15:0]   mIMOReceiverUnit_14_shift_q_6;
  wire       [15:0]   mIMOReceiverUnit_14_shift_q_7;
  wire       [15:0]   mIMOReceiverUnit_15_shift_i_0;
  wire       [15:0]   mIMOReceiverUnit_15_shift_i_1;
  wire       [15:0]   mIMOReceiverUnit_15_shift_i_2;
  wire       [15:0]   mIMOReceiverUnit_15_shift_i_3;
  wire       [15:0]   mIMOReceiverUnit_15_shift_i_4;
  wire       [15:0]   mIMOReceiverUnit_15_shift_i_5;
  wire       [15:0]   mIMOReceiverUnit_15_shift_i_6;
  wire       [15:0]   mIMOReceiverUnit_15_shift_i_7;
  wire       [15:0]   mIMOReceiverUnit_15_shift_q_0;
  wire       [15:0]   mIMOReceiverUnit_15_shift_q_1;
  wire       [15:0]   mIMOReceiverUnit_15_shift_q_2;
  wire       [15:0]   mIMOReceiverUnit_15_shift_q_3;
  wire       [15:0]   mIMOReceiverUnit_15_shift_q_4;
  wire       [15:0]   mIMOReceiverUnit_15_shift_q_5;
  wire       [15:0]   mIMOReceiverUnit_15_shift_q_6;
  wire       [15:0]   mIMOReceiverUnit_15_shift_q_7;
  wire                mIMOReceiverUnit_8_base_sub_iq_valid;
  wire       [31:0]   mIMOReceiverUnit_8_base_sub_iq_payload_cha_i;
  wire       [31:0]   mIMOReceiverUnit_8_base_sub_iq_payload_cha_q;
  wire                mIMOReceiverUnit_9_base_sub_iq_valid;
  wire       [31:0]   mIMOReceiverUnit_9_base_sub_iq_payload_cha_i;
  wire       [31:0]   mIMOReceiverUnit_9_base_sub_iq_payload_cha_q;
  wire                mIMOReceiverUnit_10_base_sub_iq_valid;
  wire       [31:0]   mIMOReceiverUnit_10_base_sub_iq_payload_cha_i;
  wire       [31:0]   mIMOReceiverUnit_10_base_sub_iq_payload_cha_q;
  wire                mIMOReceiverUnit_11_base_sub_iq_valid;
  wire       [31:0]   mIMOReceiverUnit_11_base_sub_iq_payload_cha_i;
  wire       [31:0]   mIMOReceiverUnit_11_base_sub_iq_payload_cha_q;
  wire                mIMOReceiverUnit_12_base_sub_iq_valid;
  wire       [31:0]   mIMOReceiverUnit_12_base_sub_iq_payload_cha_i;
  wire       [31:0]   mIMOReceiverUnit_12_base_sub_iq_payload_cha_q;
  wire                mIMOReceiverUnit_13_base_sub_iq_valid;
  wire       [31:0]   mIMOReceiverUnit_13_base_sub_iq_payload_cha_i;
  wire       [31:0]   mIMOReceiverUnit_13_base_sub_iq_payload_cha_q;
  wire                mIMOReceiverUnit_14_base_sub_iq_valid;
  wire       [31:0]   mIMOReceiverUnit_14_base_sub_iq_payload_cha_i;
  wire       [31:0]   mIMOReceiverUnit_14_base_sub_iq_payload_cha_q;
  wire                mIMOReceiverUnit_15_base_sub_iq_valid;
  wire       [31:0]   mIMOReceiverUnit_15_base_sub_iq_payload_cha_i;
  wire       [31:0]   mIMOReceiverUnit_15_base_sub_iq_payload_cha_q;
  reg        [15:0]   _zz_shift_i_0;
  wire       [5:0]    _zz_shift_i_0_1;
  reg        [15:0]   _zz_shift_q_0;
  wire       [5:0]    _zz_shift_q_0_1;
  reg        [15:0]   _zz_shift_i_1;
  wire       [5:0]    _zz_shift_i_1_1;
  reg        [15:0]   _zz_shift_q_1;
  wire       [5:0]    _zz_shift_q_1_1;
  reg        [15:0]   _zz_shift_i_2;
  wire       [5:0]    _zz_shift_i_2_1;
  reg        [15:0]   _zz_shift_q_2;
  wire       [5:0]    _zz_shift_q_2_1;
  reg        [15:0]   _zz_shift_i_3;
  wire       [5:0]    _zz_shift_i_3_1;
  reg        [15:0]   _zz_shift_q_3;
  wire       [5:0]    _zz_shift_q_3_1;
  reg        [15:0]   _zz_shift_i_4;
  wire       [5:0]    _zz_shift_i_4_1;
  reg        [15:0]   _zz_shift_q_4;
  wire       [5:0]    _zz_shift_q_4_1;
  reg        [15:0]   _zz_shift_i_5;
  wire       [5:0]    _zz_shift_i_5_1;
  reg        [15:0]   _zz_shift_q_5;
  wire       [5:0]    _zz_shift_q_5_1;
  reg        [15:0]   _zz_shift_i_6;
  wire       [5:0]    _zz_shift_i_6_1;
  reg        [15:0]   _zz_shift_q_6;
  wire       [5:0]    _zz_shift_q_6_1;
  reg        [15:0]   _zz_shift_i_7;
  wire       [5:0]    _zz_shift_i_7_1;
  reg        [15:0]   _zz_shift_q_7;
  wire       [5:0]    _zz_shift_q_7_1;
  reg        [15:0]   _zz_shift_i_0_2;
  wire       [5:0]    _zz_shift_i_0_3;
  reg        [15:0]   _zz_shift_q_0_2;
  wire       [5:0]    _zz_shift_q_0_3;
  reg        [15:0]   _zz_shift_i_1_2;
  wire       [5:0]    _zz_shift_i_1_3;
  reg        [15:0]   _zz_shift_q_1_2;
  wire       [5:0]    _zz_shift_q_1_3;
  reg        [15:0]   _zz_shift_i_2_2;
  wire       [5:0]    _zz_shift_i_2_3;
  reg        [15:0]   _zz_shift_q_2_2;
  wire       [5:0]    _zz_shift_q_2_3;
  reg        [15:0]   _zz_shift_i_3_2;
  wire       [5:0]    _zz_shift_i_3_3;
  reg        [15:0]   _zz_shift_q_3_2;
  wire       [5:0]    _zz_shift_q_3_3;
  reg        [15:0]   _zz_shift_i_4_2;
  wire       [5:0]    _zz_shift_i_4_3;
  reg        [15:0]   _zz_shift_q_4_2;
  wire       [5:0]    _zz_shift_q_4_3;
  reg        [15:0]   _zz_shift_i_5_2;
  wire       [5:0]    _zz_shift_i_5_3;
  reg        [15:0]   _zz_shift_q_5_2;
  wire       [5:0]    _zz_shift_q_5_3;
  reg        [15:0]   _zz_shift_i_6_2;
  wire       [5:0]    _zz_shift_i_6_3;
  reg        [15:0]   _zz_shift_q_6_2;
  wire       [5:0]    _zz_shift_q_6_3;
  reg        [15:0]   _zz_shift_i_7_2;
  wire       [5:0]    _zz_shift_i_7_3;
  reg        [15:0]   _zz_shift_q_7_2;
  wire       [5:0]    _zz_shift_q_7_3;
  reg        [15:0]   _zz_shift_i_0_4;
  wire       [5:0]    _zz_shift_i_0_5;
  reg        [15:0]   _zz_shift_q_0_4;
  wire       [5:0]    _zz_shift_q_0_5;
  reg        [15:0]   _zz_shift_i_1_4;
  wire       [5:0]    _zz_shift_i_1_5;
  reg        [15:0]   _zz_shift_q_1_4;
  wire       [5:0]    _zz_shift_q_1_5;
  reg        [15:0]   _zz_shift_i_2_4;
  wire       [5:0]    _zz_shift_i_2_5;
  reg        [15:0]   _zz_shift_q_2_4;
  wire       [5:0]    _zz_shift_q_2_5;
  reg        [15:0]   _zz_shift_i_3_4;
  wire       [5:0]    _zz_shift_i_3_5;
  reg        [15:0]   _zz_shift_q_3_4;
  wire       [5:0]    _zz_shift_q_3_5;
  reg        [15:0]   _zz_shift_i_4_4;
  wire       [5:0]    _zz_shift_i_4_5;
  reg        [15:0]   _zz_shift_q_4_4;
  wire       [5:0]    _zz_shift_q_4_5;
  reg        [15:0]   _zz_shift_i_5_4;
  wire       [5:0]    _zz_shift_i_5_5;
  reg        [15:0]   _zz_shift_q_5_4;
  wire       [5:0]    _zz_shift_q_5_5;
  reg        [15:0]   _zz_shift_i_6_4;
  wire       [5:0]    _zz_shift_i_6_5;
  reg        [15:0]   _zz_shift_q_6_4;
  wire       [5:0]    _zz_shift_q_6_5;
  reg        [15:0]   _zz_shift_i_7_4;
  wire       [5:0]    _zz_shift_i_7_5;
  reg        [15:0]   _zz_shift_q_7_4;
  wire       [5:0]    _zz_shift_q_7_5;
  reg        [15:0]   _zz_shift_i_0_6;
  wire       [5:0]    _zz_shift_i_0_7;
  reg        [15:0]   _zz_shift_q_0_6;
  wire       [5:0]    _zz_shift_q_0_7;
  reg        [15:0]   _zz_shift_i_1_6;
  wire       [5:0]    _zz_shift_i_1_7;
  reg        [15:0]   _zz_shift_q_1_6;
  wire       [5:0]    _zz_shift_q_1_7;
  reg        [15:0]   _zz_shift_i_2_6;
  wire       [5:0]    _zz_shift_i_2_7;
  reg        [15:0]   _zz_shift_q_2_6;
  wire       [5:0]    _zz_shift_q_2_7;
  reg        [15:0]   _zz_shift_i_3_6;
  wire       [5:0]    _zz_shift_i_3_7;
  reg        [15:0]   _zz_shift_q_3_6;
  wire       [5:0]    _zz_shift_q_3_7;
  reg        [15:0]   _zz_shift_i_4_6;
  wire       [5:0]    _zz_shift_i_4_7;
  reg        [15:0]   _zz_shift_q_4_6;
  wire       [5:0]    _zz_shift_q_4_7;
  reg        [15:0]   _zz_shift_i_5_6;
  wire       [5:0]    _zz_shift_i_5_7;
  reg        [15:0]   _zz_shift_q_5_6;
  wire       [5:0]    _zz_shift_q_5_7;
  reg        [15:0]   _zz_shift_i_6_6;
  wire       [5:0]    _zz_shift_i_6_7;
  reg        [15:0]   _zz_shift_q_6_6;
  wire       [5:0]    _zz_shift_q_6_7;
  reg        [15:0]   _zz_shift_i_7_6;
  wire       [5:0]    _zz_shift_i_7_7;
  reg        [15:0]   _zz_shift_q_7_6;
  wire       [5:0]    _zz_shift_q_7_7;
  reg        [15:0]   _zz_shift_i_0_8;
  wire       [5:0]    _zz_shift_i_0_9;
  reg        [15:0]   _zz_shift_q_0_8;
  wire       [5:0]    _zz_shift_q_0_9;
  reg        [15:0]   _zz_shift_i_1_8;
  wire       [5:0]    _zz_shift_i_1_9;
  reg        [15:0]   _zz_shift_q_1_8;
  wire       [5:0]    _zz_shift_q_1_9;
  reg        [15:0]   _zz_shift_i_2_8;
  wire       [5:0]    _zz_shift_i_2_9;
  reg        [15:0]   _zz_shift_q_2_8;
  wire       [5:0]    _zz_shift_q_2_9;
  reg        [15:0]   _zz_shift_i_3_8;
  wire       [5:0]    _zz_shift_i_3_9;
  reg        [15:0]   _zz_shift_q_3_8;
  wire       [5:0]    _zz_shift_q_3_9;
  reg        [15:0]   _zz_shift_i_4_8;
  wire       [5:0]    _zz_shift_i_4_9;
  reg        [15:0]   _zz_shift_q_4_8;
  wire       [5:0]    _zz_shift_q_4_9;
  reg        [15:0]   _zz_shift_i_5_8;
  wire       [5:0]    _zz_shift_i_5_9;
  reg        [15:0]   _zz_shift_q_5_8;
  wire       [5:0]    _zz_shift_q_5_9;
  reg        [15:0]   _zz_shift_i_6_8;
  wire       [5:0]    _zz_shift_i_6_9;
  reg        [15:0]   _zz_shift_q_6_8;
  wire       [5:0]    _zz_shift_q_6_9;
  reg        [15:0]   _zz_shift_i_7_8;
  wire       [5:0]    _zz_shift_i_7_9;
  reg        [15:0]   _zz_shift_q_7_8;
  wire       [5:0]    _zz_shift_q_7_9;
  reg        [15:0]   _zz_shift_i_0_10;
  wire       [5:0]    _zz_shift_i_0_11;
  reg        [15:0]   _zz_shift_q_0_10;
  wire       [5:0]    _zz_shift_q_0_11;
  reg        [15:0]   _zz_shift_i_1_10;
  wire       [5:0]    _zz_shift_i_1_11;
  reg        [15:0]   _zz_shift_q_1_10;
  wire       [5:0]    _zz_shift_q_1_11;
  reg        [15:0]   _zz_shift_i_2_10;
  wire       [5:0]    _zz_shift_i_2_11;
  reg        [15:0]   _zz_shift_q_2_10;
  wire       [5:0]    _zz_shift_q_2_11;
  reg        [15:0]   _zz_shift_i_3_10;
  wire       [5:0]    _zz_shift_i_3_11;
  reg        [15:0]   _zz_shift_q_3_10;
  wire       [5:0]    _zz_shift_q_3_11;
  reg        [15:0]   _zz_shift_i_4_10;
  wire       [5:0]    _zz_shift_i_4_11;
  reg        [15:0]   _zz_shift_q_4_10;
  wire       [5:0]    _zz_shift_q_4_11;
  reg        [15:0]   _zz_shift_i_5_10;
  wire       [5:0]    _zz_shift_i_5_11;
  reg        [15:0]   _zz_shift_q_5_10;
  wire       [5:0]    _zz_shift_q_5_11;
  reg        [15:0]   _zz_shift_i_6_10;
  wire       [5:0]    _zz_shift_i_6_11;
  reg        [15:0]   _zz_shift_q_6_10;
  wire       [5:0]    _zz_shift_q_6_11;
  reg        [15:0]   _zz_shift_i_7_10;
  wire       [5:0]    _zz_shift_i_7_11;
  reg        [15:0]   _zz_shift_q_7_10;
  wire       [5:0]    _zz_shift_q_7_11;
  reg        [15:0]   _zz_shift_i_0_12;
  wire       [5:0]    _zz_shift_i_0_13;
  reg        [15:0]   _zz_shift_q_0_12;
  wire       [5:0]    _zz_shift_q_0_13;
  reg        [15:0]   _zz_shift_i_1_12;
  wire       [5:0]    _zz_shift_i_1_13;
  reg        [15:0]   _zz_shift_q_1_12;
  wire       [5:0]    _zz_shift_q_1_13;
  reg        [15:0]   _zz_shift_i_2_12;
  wire       [5:0]    _zz_shift_i_2_13;
  reg        [15:0]   _zz_shift_q_2_12;
  wire       [5:0]    _zz_shift_q_2_13;
  reg        [15:0]   _zz_shift_i_3_12;
  wire       [5:0]    _zz_shift_i_3_13;
  reg        [15:0]   _zz_shift_q_3_12;
  wire       [5:0]    _zz_shift_q_3_13;
  reg        [15:0]   _zz_shift_i_4_12;
  wire       [5:0]    _zz_shift_i_4_13;
  reg        [15:0]   _zz_shift_q_4_12;
  wire       [5:0]    _zz_shift_q_4_13;
  reg        [15:0]   _zz_shift_i_5_12;
  wire       [5:0]    _zz_shift_i_5_13;
  reg        [15:0]   _zz_shift_q_5_12;
  wire       [5:0]    _zz_shift_q_5_13;
  reg        [15:0]   _zz_shift_i_6_12;
  wire       [5:0]    _zz_shift_i_6_13;
  reg        [15:0]   _zz_shift_q_6_12;
  wire       [5:0]    _zz_shift_q_6_13;
  reg        [15:0]   _zz_shift_i_7_12;
  wire       [5:0]    _zz_shift_i_7_13;
  reg        [15:0]   _zz_shift_q_7_12;
  wire       [5:0]    _zz_shift_q_7_13;
  reg        [15:0]   _zz_shift_i_0_14;
  wire       [5:0]    _zz_shift_i_0_15;
  reg        [15:0]   _zz_shift_q_0_14;
  wire       [5:0]    _zz_shift_q_0_15;
  reg        [15:0]   _zz_shift_i_1_14;
  wire       [5:0]    _zz_shift_i_1_15;
  reg        [15:0]   _zz_shift_q_1_14;
  wire       [5:0]    _zz_shift_q_1_15;
  reg        [15:0]   _zz_shift_i_2_14;
  wire       [5:0]    _zz_shift_i_2_15;
  reg        [15:0]   _zz_shift_q_2_14;
  wire       [5:0]    _zz_shift_q_2_15;
  reg        [15:0]   _zz_shift_i_3_14;
  wire       [5:0]    _zz_shift_i_3_15;
  reg        [15:0]   _zz_shift_q_3_14;
  wire       [5:0]    _zz_shift_q_3_15;
  reg        [15:0]   _zz_shift_i_4_14;
  wire       [5:0]    _zz_shift_i_4_15;
  reg        [15:0]   _zz_shift_q_4_14;
  wire       [5:0]    _zz_shift_q_4_15;
  reg        [15:0]   _zz_shift_i_5_14;
  wire       [5:0]    _zz_shift_i_5_15;
  reg        [15:0]   _zz_shift_q_5_14;
  wire       [5:0]    _zz_shift_q_5_15;
  reg        [15:0]   _zz_shift_i_6_14;
  wire       [5:0]    _zz_shift_i_6_15;
  reg        [15:0]   _zz_shift_q_6_14;
  wire       [5:0]    _zz_shift_q_6_15;
  reg        [15:0]   _zz_shift_i_7_14;
  wire       [5:0]    _zz_shift_i_7_15;
  reg        [15:0]   _zz_shift_q_7_14;
  wire       [5:0]    _zz_shift_q_7_15;
  reg        [15:0]   shift_i_map_0;
  reg        [15:0]   shift_i_map_1;
  reg        [15:0]   shift_i_map_2;
  reg        [15:0]   shift_i_map_3;
  reg        [15:0]   shift_i_map_4;
  reg        [15:0]   shift_i_map_5;
  reg        [15:0]   shift_i_map_6;
  reg        [15:0]   shift_i_map_7;
  reg        [15:0]   shift_i_map_8;
  reg        [15:0]   shift_i_map_9;
  reg        [15:0]   shift_i_map_10;
  reg        [15:0]   shift_i_map_11;
  reg        [15:0]   shift_i_map_12;
  reg        [15:0]   shift_i_map_13;
  reg        [15:0]   shift_i_map_14;
  reg        [15:0]   shift_i_map_15;
  reg        [15:0]   shift_i_map_16;
  reg        [15:0]   shift_i_map_17;
  reg        [15:0]   shift_i_map_18;
  reg        [15:0]   shift_i_map_19;
  reg        [15:0]   shift_i_map_20;
  reg        [15:0]   shift_i_map_21;
  reg        [15:0]   shift_i_map_22;
  reg        [15:0]   shift_i_map_23;
  reg        [15:0]   shift_i_map_24;
  reg        [15:0]   shift_i_map_25;
  reg        [15:0]   shift_i_map_26;
  reg        [15:0]   shift_i_map_27;
  reg        [15:0]   shift_i_map_28;
  reg        [15:0]   shift_i_map_29;
  reg        [15:0]   shift_i_map_30;
  reg        [15:0]   shift_i_map_31;
  reg        [15:0]   shift_i_map_32;
  reg        [15:0]   shift_i_map_33;
  reg        [15:0]   shift_i_map_34;
  reg        [15:0]   shift_i_map_35;
  reg        [15:0]   shift_i_map_36;
  reg        [15:0]   shift_i_map_37;
  reg        [15:0]   shift_i_map_38;
  reg        [15:0]   shift_i_map_39;
  reg        [15:0]   shift_i_map_40;
  reg        [15:0]   shift_i_map_41;
  reg        [15:0]   shift_i_map_42;
  reg        [15:0]   shift_i_map_43;
  reg        [15:0]   shift_i_map_44;
  reg        [15:0]   shift_i_map_45;
  reg        [15:0]   shift_i_map_46;
  reg        [15:0]   shift_i_map_47;
  reg        [15:0]   shift_i_map_48;
  reg        [15:0]   shift_i_map_49;
  reg        [15:0]   shift_i_map_50;
  reg        [15:0]   shift_i_map_51;
  reg        [15:0]   shift_i_map_52;
  reg        [15:0]   shift_i_map_53;
  reg        [15:0]   shift_i_map_54;
  reg        [15:0]   shift_i_map_55;
  reg        [15:0]   shift_i_map_56;
  reg        [15:0]   shift_i_map_57;
  reg        [15:0]   shift_i_map_58;
  reg        [15:0]   shift_i_map_59;
  reg        [15:0]   shift_i_map_60;
  reg        [15:0]   shift_i_map_61;
  reg        [15:0]   shift_i_map_62;
  reg        [15:0]   shift_i_map_63;
  reg        [15:0]   shift_q_map_0;
  reg        [15:0]   shift_q_map_1;
  reg        [15:0]   shift_q_map_2;
  reg        [15:0]   shift_q_map_3;
  reg        [15:0]   shift_q_map_4;
  reg        [15:0]   shift_q_map_5;
  reg        [15:0]   shift_q_map_6;
  reg        [15:0]   shift_q_map_7;
  reg        [15:0]   shift_q_map_8;
  reg        [15:0]   shift_q_map_9;
  reg        [15:0]   shift_q_map_10;
  reg        [15:0]   shift_q_map_11;
  reg        [15:0]   shift_q_map_12;
  reg        [15:0]   shift_q_map_13;
  reg        [15:0]   shift_q_map_14;
  reg        [15:0]   shift_q_map_15;
  reg        [15:0]   shift_q_map_16;
  reg        [15:0]   shift_q_map_17;
  reg        [15:0]   shift_q_map_18;
  reg        [15:0]   shift_q_map_19;
  reg        [15:0]   shift_q_map_20;
  reg        [15:0]   shift_q_map_21;
  reg        [15:0]   shift_q_map_22;
  reg        [15:0]   shift_q_map_23;
  reg        [15:0]   shift_q_map_24;
  reg        [15:0]   shift_q_map_25;
  reg        [15:0]   shift_q_map_26;
  reg        [15:0]   shift_q_map_27;
  reg        [15:0]   shift_q_map_28;
  reg        [15:0]   shift_q_map_29;
  reg        [15:0]   shift_q_map_30;
  reg        [15:0]   shift_q_map_31;
  reg        [15:0]   shift_q_map_32;
  reg        [15:0]   shift_q_map_33;
  reg        [15:0]   shift_q_map_34;
  reg        [15:0]   shift_q_map_35;
  reg        [15:0]   shift_q_map_36;
  reg        [15:0]   shift_q_map_37;
  reg        [15:0]   shift_q_map_38;
  reg        [15:0]   shift_q_map_39;
  reg        [15:0]   shift_q_map_40;
  reg        [15:0]   shift_q_map_41;
  reg        [15:0]   shift_q_map_42;
  reg        [15:0]   shift_q_map_43;
  reg        [15:0]   shift_q_map_44;
  reg        [15:0]   shift_q_map_45;
  reg        [15:0]   shift_q_map_46;
  reg        [15:0]   shift_q_map_47;
  reg        [15:0]   shift_q_map_48;
  reg        [15:0]   shift_q_map_49;
  reg        [15:0]   shift_q_map_50;
  reg        [15:0]   shift_q_map_51;
  reg        [15:0]   shift_q_map_52;
  reg        [15:0]   shift_q_map_53;
  reg        [15:0]   shift_q_map_54;
  reg        [15:0]   shift_q_map_55;
  reg        [15:0]   shift_q_map_56;
  reg        [15:0]   shift_q_map_57;
  reg        [15:0]   shift_q_map_58;
  reg        [15:0]   shift_q_map_59;
  reg        [15:0]   shift_q_map_60;
  reg        [15:0]   shift_q_map_61;
  reg        [15:0]   shift_q_map_62;
  reg        [15:0]   shift_q_map_63;
  wire       [63:0]   _zz_1;
  wire       [63:0]   _zz_2;
  wire                base_sub_valid_vec_0;
  wire                base_sub_valid_vec_1;
  wire                base_sub_valid_vec_2;
  wire                base_sub_valid_vec_3;
  wire                base_sub_valid_vec_4;
  wire                base_sub_valid_vec_5;
  wire                base_sub_valid_vec_6;
  wire                base_sub_valid_vec_7;

  assign _zz_shift_i_0_1 = 6'h0;
  assign _zz_shift_q_0_1 = 6'h0;
  assign _zz_shift_i_1_1 = 6'h01;
  assign _zz_shift_q_1_1 = 6'h01;
  assign _zz_shift_i_2_1 = 6'h02;
  assign _zz_shift_q_2_1 = 6'h02;
  assign _zz_shift_i_3_1 = 6'h03;
  assign _zz_shift_q_3_1 = 6'h03;
  assign _zz_shift_i_4_1 = 6'h04;
  assign _zz_shift_q_4_1 = 6'h04;
  assign _zz_shift_i_5_1 = 6'h05;
  assign _zz_shift_q_5_1 = 6'h05;
  assign _zz_shift_i_6_1 = 6'h06;
  assign _zz_shift_q_6_1 = 6'h06;
  assign _zz_shift_i_7_1 = 6'h07;
  assign _zz_shift_q_7_1 = 6'h07;
  assign _zz_shift_i_0_3 = 6'h08;
  assign _zz_shift_q_0_3 = 6'h08;
  assign _zz_shift_i_1_3 = 6'h09;
  assign _zz_shift_q_1_3 = 6'h09;
  assign _zz_shift_i_2_3 = 6'h0a;
  assign _zz_shift_q_2_3 = 6'h0a;
  assign _zz_shift_i_3_3 = 6'h0b;
  assign _zz_shift_q_3_3 = 6'h0b;
  assign _zz_shift_i_4_3 = 6'h0c;
  assign _zz_shift_q_4_3 = 6'h0c;
  assign _zz_shift_i_5_3 = 6'h0d;
  assign _zz_shift_q_5_3 = 6'h0d;
  assign _zz_shift_i_6_3 = 6'h0e;
  assign _zz_shift_q_6_3 = 6'h0e;
  assign _zz_shift_i_7_3 = 6'h0f;
  assign _zz_shift_q_7_3 = 6'h0f;
  assign _zz_shift_i_0_5 = 6'h10;
  assign _zz_shift_q_0_5 = 6'h10;
  assign _zz_shift_i_1_5 = 6'h11;
  assign _zz_shift_q_1_5 = 6'h11;
  assign _zz_shift_i_2_5 = 6'h12;
  assign _zz_shift_q_2_5 = 6'h12;
  assign _zz_shift_i_3_5 = 6'h13;
  assign _zz_shift_q_3_5 = 6'h13;
  assign _zz_shift_i_4_5 = 6'h14;
  assign _zz_shift_q_4_5 = 6'h14;
  assign _zz_shift_i_5_5 = 6'h15;
  assign _zz_shift_q_5_5 = 6'h15;
  assign _zz_shift_i_6_5 = 6'h16;
  assign _zz_shift_q_6_5 = 6'h16;
  assign _zz_shift_i_7_5 = 6'h17;
  assign _zz_shift_q_7_5 = 6'h17;
  assign _zz_shift_i_0_7 = 6'h18;
  assign _zz_shift_q_0_7 = 6'h18;
  assign _zz_shift_i_1_7 = 6'h19;
  assign _zz_shift_q_1_7 = 6'h19;
  assign _zz_shift_i_2_7 = 6'h1a;
  assign _zz_shift_q_2_7 = 6'h1a;
  assign _zz_shift_i_3_7 = 6'h1b;
  assign _zz_shift_q_3_7 = 6'h1b;
  assign _zz_shift_i_4_7 = 6'h1c;
  assign _zz_shift_q_4_7 = 6'h1c;
  assign _zz_shift_i_5_7 = 6'h1d;
  assign _zz_shift_q_5_7 = 6'h1d;
  assign _zz_shift_i_6_7 = 6'h1e;
  assign _zz_shift_q_6_7 = 6'h1e;
  assign _zz_shift_i_7_7 = 6'h1f;
  assign _zz_shift_q_7_7 = 6'h1f;
  assign _zz_shift_i_0_9 = 6'h20;
  assign _zz_shift_q_0_9 = 6'h20;
  assign _zz_shift_i_1_9 = 6'h21;
  assign _zz_shift_q_1_9 = 6'h21;
  assign _zz_shift_i_2_9 = 6'h22;
  assign _zz_shift_q_2_9 = 6'h22;
  assign _zz_shift_i_3_9 = 6'h23;
  assign _zz_shift_q_3_9 = 6'h23;
  assign _zz_shift_i_4_9 = 6'h24;
  assign _zz_shift_q_4_9 = 6'h24;
  assign _zz_shift_i_5_9 = 6'h25;
  assign _zz_shift_q_5_9 = 6'h25;
  assign _zz_shift_i_6_9 = 6'h26;
  assign _zz_shift_q_6_9 = 6'h26;
  assign _zz_shift_i_7_9 = 6'h27;
  assign _zz_shift_q_7_9 = 6'h27;
  assign _zz_shift_i_0_11 = 6'h28;
  assign _zz_shift_q_0_11 = 6'h28;
  assign _zz_shift_i_1_11 = 6'h29;
  assign _zz_shift_q_1_11 = 6'h29;
  assign _zz_shift_i_2_11 = 6'h2a;
  assign _zz_shift_q_2_11 = 6'h2a;
  assign _zz_shift_i_3_11 = 6'h2b;
  assign _zz_shift_q_3_11 = 6'h2b;
  assign _zz_shift_i_4_11 = 6'h2c;
  assign _zz_shift_q_4_11 = 6'h2c;
  assign _zz_shift_i_5_11 = 6'h2d;
  assign _zz_shift_q_5_11 = 6'h2d;
  assign _zz_shift_i_6_11 = 6'h2e;
  assign _zz_shift_q_6_11 = 6'h2e;
  assign _zz_shift_i_7_11 = 6'h2f;
  assign _zz_shift_q_7_11 = 6'h2f;
  assign _zz_shift_i_0_13 = 6'h30;
  assign _zz_shift_q_0_13 = 6'h30;
  assign _zz_shift_i_1_13 = 6'h31;
  assign _zz_shift_q_1_13 = 6'h31;
  assign _zz_shift_i_2_13 = 6'h32;
  assign _zz_shift_q_2_13 = 6'h32;
  assign _zz_shift_i_3_13 = 6'h33;
  assign _zz_shift_q_3_13 = 6'h33;
  assign _zz_shift_i_4_13 = 6'h34;
  assign _zz_shift_q_4_13 = 6'h34;
  assign _zz_shift_i_5_13 = 6'h35;
  assign _zz_shift_q_5_13 = 6'h35;
  assign _zz_shift_i_6_13 = 6'h36;
  assign _zz_shift_q_6_13 = 6'h36;
  assign _zz_shift_i_7_13 = 6'h37;
  assign _zz_shift_q_7_13 = 6'h37;
  assign _zz_shift_i_0_15 = 6'h38;
  assign _zz_shift_q_0_15 = 6'h38;
  assign _zz_shift_i_1_15 = 6'h39;
  assign _zz_shift_q_1_15 = 6'h39;
  assign _zz_shift_i_2_15 = 6'h3a;
  assign _zz_shift_q_2_15 = 6'h3a;
  assign _zz_shift_i_3_15 = 6'h3b;
  assign _zz_shift_q_3_15 = 6'h3b;
  assign _zz_shift_i_4_15 = 6'h3c;
  assign _zz_shift_q_4_15 = 6'h3c;
  assign _zz_shift_i_5_15 = 6'h3d;
  assign _zz_shift_q_5_15 = 6'h3d;
  assign _zz_shift_i_6_15 = 6'h3e;
  assign _zz_shift_q_6_15 = 6'h3e;
  assign _zz_shift_i_7_15 = 6'h3f;
  assign _zz_shift_q_7_15 = 6'h3f;
  MIMOReceiverUnit mIMOReceiverUnit_8 (
    .shift_i_0                 (mIMOReceiverUnit_8_shift_i_0[15:0]                ), //i
    .shift_i_1                 (mIMOReceiverUnit_8_shift_i_1[15:0]                ), //i
    .shift_i_2                 (mIMOReceiverUnit_8_shift_i_2[15:0]                ), //i
    .shift_i_3                 (mIMOReceiverUnit_8_shift_i_3[15:0]                ), //i
    .shift_i_4                 (mIMOReceiverUnit_8_shift_i_4[15:0]                ), //i
    .shift_i_5                 (mIMOReceiverUnit_8_shift_i_5[15:0]                ), //i
    .shift_i_6                 (mIMOReceiverUnit_8_shift_i_6[15:0]                ), //i
    .shift_i_7                 (mIMOReceiverUnit_8_shift_i_7[15:0]                ), //i
    .shift_q_0                 (mIMOReceiverUnit_8_shift_q_0[15:0]                ), //i
    .shift_q_1                 (mIMOReceiverUnit_8_shift_q_1[15:0]                ), //i
    .shift_q_2                 (mIMOReceiverUnit_8_shift_q_2[15:0]                ), //i
    .shift_q_3                 (mIMOReceiverUnit_8_shift_q_3[15:0]                ), //i
    .shift_q_4                 (mIMOReceiverUnit_8_shift_q_4[15:0]                ), //i
    .shift_q_5                 (mIMOReceiverUnit_8_shift_q_5[15:0]                ), //i
    .shift_q_6                 (mIMOReceiverUnit_8_shift_q_6[15:0]                ), //i
    .shift_q_7                 (mIMOReceiverUnit_8_shift_q_7[15:0]                ), //i
    .mod_iq_valid              (mod_iq_valid                                      ), //i
    .mod_iq_payload_cha_i      (mod_iq_payload_cha_i[15:0]                        ), //i
    .mod_iq_payload_cha_q      (mod_iq_payload_cha_q[15:0]                        ), //i
    .base_sub_iq_valid         (mIMOReceiverUnit_8_base_sub_iq_valid              ), //o
    .base_sub_iq_payload_cha_i (mIMOReceiverUnit_8_base_sub_iq_payload_cha_i[31:0]), //o
    .base_sub_iq_payload_cha_q (mIMOReceiverUnit_8_base_sub_iq_payload_cha_q[31:0]), //o
    .rf_clk                    (rf_clk                                            ), //i
    .rf_resetn                 (rf_resetn                                         )  //i
  );
  MIMOReceiverUnit mIMOReceiverUnit_9 (
    .shift_i_0                 (mIMOReceiverUnit_9_shift_i_0[15:0]                ), //i
    .shift_i_1                 (mIMOReceiverUnit_9_shift_i_1[15:0]                ), //i
    .shift_i_2                 (mIMOReceiverUnit_9_shift_i_2[15:0]                ), //i
    .shift_i_3                 (mIMOReceiverUnit_9_shift_i_3[15:0]                ), //i
    .shift_i_4                 (mIMOReceiverUnit_9_shift_i_4[15:0]                ), //i
    .shift_i_5                 (mIMOReceiverUnit_9_shift_i_5[15:0]                ), //i
    .shift_i_6                 (mIMOReceiverUnit_9_shift_i_6[15:0]                ), //i
    .shift_i_7                 (mIMOReceiverUnit_9_shift_i_7[15:0]                ), //i
    .shift_q_0                 (mIMOReceiverUnit_9_shift_q_0[15:0]                ), //i
    .shift_q_1                 (mIMOReceiverUnit_9_shift_q_1[15:0]                ), //i
    .shift_q_2                 (mIMOReceiverUnit_9_shift_q_2[15:0]                ), //i
    .shift_q_3                 (mIMOReceiverUnit_9_shift_q_3[15:0]                ), //i
    .shift_q_4                 (mIMOReceiverUnit_9_shift_q_4[15:0]                ), //i
    .shift_q_5                 (mIMOReceiverUnit_9_shift_q_5[15:0]                ), //i
    .shift_q_6                 (mIMOReceiverUnit_9_shift_q_6[15:0]                ), //i
    .shift_q_7                 (mIMOReceiverUnit_9_shift_q_7[15:0]                ), //i
    .mod_iq_valid              (mod_iq_valid                                      ), //i
    .mod_iq_payload_cha_i      (mod_iq_payload_cha_i[15:0]                        ), //i
    .mod_iq_payload_cha_q      (mod_iq_payload_cha_q[15:0]                        ), //i
    .base_sub_iq_valid         (mIMOReceiverUnit_9_base_sub_iq_valid              ), //o
    .base_sub_iq_payload_cha_i (mIMOReceiverUnit_9_base_sub_iq_payload_cha_i[31:0]), //o
    .base_sub_iq_payload_cha_q (mIMOReceiverUnit_9_base_sub_iq_payload_cha_q[31:0]), //o
    .rf_clk                    (rf_clk                                            ), //i
    .rf_resetn                 (rf_resetn                                         )  //i
  );
  MIMOReceiverUnit mIMOReceiverUnit_10 (
    .shift_i_0                 (mIMOReceiverUnit_10_shift_i_0[15:0]                ), //i
    .shift_i_1                 (mIMOReceiverUnit_10_shift_i_1[15:0]                ), //i
    .shift_i_2                 (mIMOReceiverUnit_10_shift_i_2[15:0]                ), //i
    .shift_i_3                 (mIMOReceiverUnit_10_shift_i_3[15:0]                ), //i
    .shift_i_4                 (mIMOReceiverUnit_10_shift_i_4[15:0]                ), //i
    .shift_i_5                 (mIMOReceiverUnit_10_shift_i_5[15:0]                ), //i
    .shift_i_6                 (mIMOReceiverUnit_10_shift_i_6[15:0]                ), //i
    .shift_i_7                 (mIMOReceiverUnit_10_shift_i_7[15:0]                ), //i
    .shift_q_0                 (mIMOReceiverUnit_10_shift_q_0[15:0]                ), //i
    .shift_q_1                 (mIMOReceiverUnit_10_shift_q_1[15:0]                ), //i
    .shift_q_2                 (mIMOReceiverUnit_10_shift_q_2[15:0]                ), //i
    .shift_q_3                 (mIMOReceiverUnit_10_shift_q_3[15:0]                ), //i
    .shift_q_4                 (mIMOReceiverUnit_10_shift_q_4[15:0]                ), //i
    .shift_q_5                 (mIMOReceiverUnit_10_shift_q_5[15:0]                ), //i
    .shift_q_6                 (mIMOReceiverUnit_10_shift_q_6[15:0]                ), //i
    .shift_q_7                 (mIMOReceiverUnit_10_shift_q_7[15:0]                ), //i
    .mod_iq_valid              (mod_iq_valid                                       ), //i
    .mod_iq_payload_cha_i      (mod_iq_payload_cha_i[15:0]                         ), //i
    .mod_iq_payload_cha_q      (mod_iq_payload_cha_q[15:0]                         ), //i
    .base_sub_iq_valid         (mIMOReceiverUnit_10_base_sub_iq_valid              ), //o
    .base_sub_iq_payload_cha_i (mIMOReceiverUnit_10_base_sub_iq_payload_cha_i[31:0]), //o
    .base_sub_iq_payload_cha_q (mIMOReceiverUnit_10_base_sub_iq_payload_cha_q[31:0]), //o
    .rf_clk                    (rf_clk                                             ), //i
    .rf_resetn                 (rf_resetn                                          )  //i
  );
  MIMOReceiverUnit mIMOReceiverUnit_11 (
    .shift_i_0                 (mIMOReceiverUnit_11_shift_i_0[15:0]                ), //i
    .shift_i_1                 (mIMOReceiverUnit_11_shift_i_1[15:0]                ), //i
    .shift_i_2                 (mIMOReceiverUnit_11_shift_i_2[15:0]                ), //i
    .shift_i_3                 (mIMOReceiverUnit_11_shift_i_3[15:0]                ), //i
    .shift_i_4                 (mIMOReceiverUnit_11_shift_i_4[15:0]                ), //i
    .shift_i_5                 (mIMOReceiverUnit_11_shift_i_5[15:0]                ), //i
    .shift_i_6                 (mIMOReceiverUnit_11_shift_i_6[15:0]                ), //i
    .shift_i_7                 (mIMOReceiverUnit_11_shift_i_7[15:0]                ), //i
    .shift_q_0                 (mIMOReceiverUnit_11_shift_q_0[15:0]                ), //i
    .shift_q_1                 (mIMOReceiverUnit_11_shift_q_1[15:0]                ), //i
    .shift_q_2                 (mIMOReceiverUnit_11_shift_q_2[15:0]                ), //i
    .shift_q_3                 (mIMOReceiverUnit_11_shift_q_3[15:0]                ), //i
    .shift_q_4                 (mIMOReceiverUnit_11_shift_q_4[15:0]                ), //i
    .shift_q_5                 (mIMOReceiverUnit_11_shift_q_5[15:0]                ), //i
    .shift_q_6                 (mIMOReceiverUnit_11_shift_q_6[15:0]                ), //i
    .shift_q_7                 (mIMOReceiverUnit_11_shift_q_7[15:0]                ), //i
    .mod_iq_valid              (mod_iq_valid                                       ), //i
    .mod_iq_payload_cha_i      (mod_iq_payload_cha_i[15:0]                         ), //i
    .mod_iq_payload_cha_q      (mod_iq_payload_cha_q[15:0]                         ), //i
    .base_sub_iq_valid         (mIMOReceiverUnit_11_base_sub_iq_valid              ), //o
    .base_sub_iq_payload_cha_i (mIMOReceiverUnit_11_base_sub_iq_payload_cha_i[31:0]), //o
    .base_sub_iq_payload_cha_q (mIMOReceiverUnit_11_base_sub_iq_payload_cha_q[31:0]), //o
    .rf_clk                    (rf_clk                                             ), //i
    .rf_resetn                 (rf_resetn                                          )  //i
  );
  MIMOReceiverUnit mIMOReceiverUnit_12 (
    .shift_i_0                 (mIMOReceiverUnit_12_shift_i_0[15:0]                ), //i
    .shift_i_1                 (mIMOReceiverUnit_12_shift_i_1[15:0]                ), //i
    .shift_i_2                 (mIMOReceiverUnit_12_shift_i_2[15:0]                ), //i
    .shift_i_3                 (mIMOReceiverUnit_12_shift_i_3[15:0]                ), //i
    .shift_i_4                 (mIMOReceiverUnit_12_shift_i_4[15:0]                ), //i
    .shift_i_5                 (mIMOReceiverUnit_12_shift_i_5[15:0]                ), //i
    .shift_i_6                 (mIMOReceiverUnit_12_shift_i_6[15:0]                ), //i
    .shift_i_7                 (mIMOReceiverUnit_12_shift_i_7[15:0]                ), //i
    .shift_q_0                 (mIMOReceiverUnit_12_shift_q_0[15:0]                ), //i
    .shift_q_1                 (mIMOReceiverUnit_12_shift_q_1[15:0]                ), //i
    .shift_q_2                 (mIMOReceiverUnit_12_shift_q_2[15:0]                ), //i
    .shift_q_3                 (mIMOReceiverUnit_12_shift_q_3[15:0]                ), //i
    .shift_q_4                 (mIMOReceiverUnit_12_shift_q_4[15:0]                ), //i
    .shift_q_5                 (mIMOReceiverUnit_12_shift_q_5[15:0]                ), //i
    .shift_q_6                 (mIMOReceiverUnit_12_shift_q_6[15:0]                ), //i
    .shift_q_7                 (mIMOReceiverUnit_12_shift_q_7[15:0]                ), //i
    .mod_iq_valid              (mod_iq_valid                                       ), //i
    .mod_iq_payload_cha_i      (mod_iq_payload_cha_i[15:0]                         ), //i
    .mod_iq_payload_cha_q      (mod_iq_payload_cha_q[15:0]                         ), //i
    .base_sub_iq_valid         (mIMOReceiverUnit_12_base_sub_iq_valid              ), //o
    .base_sub_iq_payload_cha_i (mIMOReceiverUnit_12_base_sub_iq_payload_cha_i[31:0]), //o
    .base_sub_iq_payload_cha_q (mIMOReceiverUnit_12_base_sub_iq_payload_cha_q[31:0]), //o
    .rf_clk                    (rf_clk                                             ), //i
    .rf_resetn                 (rf_resetn                                          )  //i
  );
  MIMOReceiverUnit mIMOReceiverUnit_13 (
    .shift_i_0                 (mIMOReceiverUnit_13_shift_i_0[15:0]                ), //i
    .shift_i_1                 (mIMOReceiverUnit_13_shift_i_1[15:0]                ), //i
    .shift_i_2                 (mIMOReceiverUnit_13_shift_i_2[15:0]                ), //i
    .shift_i_3                 (mIMOReceiverUnit_13_shift_i_3[15:0]                ), //i
    .shift_i_4                 (mIMOReceiverUnit_13_shift_i_4[15:0]                ), //i
    .shift_i_5                 (mIMOReceiverUnit_13_shift_i_5[15:0]                ), //i
    .shift_i_6                 (mIMOReceiverUnit_13_shift_i_6[15:0]                ), //i
    .shift_i_7                 (mIMOReceiverUnit_13_shift_i_7[15:0]                ), //i
    .shift_q_0                 (mIMOReceiverUnit_13_shift_q_0[15:0]                ), //i
    .shift_q_1                 (mIMOReceiverUnit_13_shift_q_1[15:0]                ), //i
    .shift_q_2                 (mIMOReceiverUnit_13_shift_q_2[15:0]                ), //i
    .shift_q_3                 (mIMOReceiverUnit_13_shift_q_3[15:0]                ), //i
    .shift_q_4                 (mIMOReceiverUnit_13_shift_q_4[15:0]                ), //i
    .shift_q_5                 (mIMOReceiverUnit_13_shift_q_5[15:0]                ), //i
    .shift_q_6                 (mIMOReceiverUnit_13_shift_q_6[15:0]                ), //i
    .shift_q_7                 (mIMOReceiverUnit_13_shift_q_7[15:0]                ), //i
    .mod_iq_valid              (mod_iq_valid                                       ), //i
    .mod_iq_payload_cha_i      (mod_iq_payload_cha_i[15:0]                         ), //i
    .mod_iq_payload_cha_q      (mod_iq_payload_cha_q[15:0]                         ), //i
    .base_sub_iq_valid         (mIMOReceiverUnit_13_base_sub_iq_valid              ), //o
    .base_sub_iq_payload_cha_i (mIMOReceiverUnit_13_base_sub_iq_payload_cha_i[31:0]), //o
    .base_sub_iq_payload_cha_q (mIMOReceiverUnit_13_base_sub_iq_payload_cha_q[31:0]), //o
    .rf_clk                    (rf_clk                                             ), //i
    .rf_resetn                 (rf_resetn                                          )  //i
  );
  MIMOReceiverUnit mIMOReceiverUnit_14 (
    .shift_i_0                 (mIMOReceiverUnit_14_shift_i_0[15:0]                ), //i
    .shift_i_1                 (mIMOReceiverUnit_14_shift_i_1[15:0]                ), //i
    .shift_i_2                 (mIMOReceiverUnit_14_shift_i_2[15:0]                ), //i
    .shift_i_3                 (mIMOReceiverUnit_14_shift_i_3[15:0]                ), //i
    .shift_i_4                 (mIMOReceiverUnit_14_shift_i_4[15:0]                ), //i
    .shift_i_5                 (mIMOReceiverUnit_14_shift_i_5[15:0]                ), //i
    .shift_i_6                 (mIMOReceiverUnit_14_shift_i_6[15:0]                ), //i
    .shift_i_7                 (mIMOReceiverUnit_14_shift_i_7[15:0]                ), //i
    .shift_q_0                 (mIMOReceiverUnit_14_shift_q_0[15:0]                ), //i
    .shift_q_1                 (mIMOReceiverUnit_14_shift_q_1[15:0]                ), //i
    .shift_q_2                 (mIMOReceiverUnit_14_shift_q_2[15:0]                ), //i
    .shift_q_3                 (mIMOReceiverUnit_14_shift_q_3[15:0]                ), //i
    .shift_q_4                 (mIMOReceiverUnit_14_shift_q_4[15:0]                ), //i
    .shift_q_5                 (mIMOReceiverUnit_14_shift_q_5[15:0]                ), //i
    .shift_q_6                 (mIMOReceiverUnit_14_shift_q_6[15:0]                ), //i
    .shift_q_7                 (mIMOReceiverUnit_14_shift_q_7[15:0]                ), //i
    .mod_iq_valid              (mod_iq_valid                                       ), //i
    .mod_iq_payload_cha_i      (mod_iq_payload_cha_i[15:0]                         ), //i
    .mod_iq_payload_cha_q      (mod_iq_payload_cha_q[15:0]                         ), //i
    .base_sub_iq_valid         (mIMOReceiverUnit_14_base_sub_iq_valid              ), //o
    .base_sub_iq_payload_cha_i (mIMOReceiverUnit_14_base_sub_iq_payload_cha_i[31:0]), //o
    .base_sub_iq_payload_cha_q (mIMOReceiverUnit_14_base_sub_iq_payload_cha_q[31:0]), //o
    .rf_clk                    (rf_clk                                             ), //i
    .rf_resetn                 (rf_resetn                                          )  //i
  );
  MIMOReceiverUnit mIMOReceiverUnit_15 (
    .shift_i_0                 (mIMOReceiverUnit_15_shift_i_0[15:0]                ), //i
    .shift_i_1                 (mIMOReceiverUnit_15_shift_i_1[15:0]                ), //i
    .shift_i_2                 (mIMOReceiverUnit_15_shift_i_2[15:0]                ), //i
    .shift_i_3                 (mIMOReceiverUnit_15_shift_i_3[15:0]                ), //i
    .shift_i_4                 (mIMOReceiverUnit_15_shift_i_4[15:0]                ), //i
    .shift_i_5                 (mIMOReceiverUnit_15_shift_i_5[15:0]                ), //i
    .shift_i_6                 (mIMOReceiverUnit_15_shift_i_6[15:0]                ), //i
    .shift_i_7                 (mIMOReceiverUnit_15_shift_i_7[15:0]                ), //i
    .shift_q_0                 (mIMOReceiverUnit_15_shift_q_0[15:0]                ), //i
    .shift_q_1                 (mIMOReceiverUnit_15_shift_q_1[15:0]                ), //i
    .shift_q_2                 (mIMOReceiverUnit_15_shift_q_2[15:0]                ), //i
    .shift_q_3                 (mIMOReceiverUnit_15_shift_q_3[15:0]                ), //i
    .shift_q_4                 (mIMOReceiverUnit_15_shift_q_4[15:0]                ), //i
    .shift_q_5                 (mIMOReceiverUnit_15_shift_q_5[15:0]                ), //i
    .shift_q_6                 (mIMOReceiverUnit_15_shift_q_6[15:0]                ), //i
    .shift_q_7                 (mIMOReceiverUnit_15_shift_q_7[15:0]                ), //i
    .mod_iq_valid              (mod_iq_valid                                       ), //i
    .mod_iq_payload_cha_i      (mod_iq_payload_cha_i[15:0]                         ), //i
    .mod_iq_payload_cha_q      (mod_iq_payload_cha_q[15:0]                         ), //i
    .base_sub_iq_valid         (mIMOReceiverUnit_15_base_sub_iq_valid              ), //o
    .base_sub_iq_payload_cha_i (mIMOReceiverUnit_15_base_sub_iq_payload_cha_i[31:0]), //o
    .base_sub_iq_payload_cha_q (mIMOReceiverUnit_15_base_sub_iq_payload_cha_q[31:0]), //o
    .rf_clk                    (rf_clk                                             ), //i
    .rf_resetn                 (rf_resetn                                          )  //i
  );
  always @(*) begin
    case(_zz_shift_i_0_1)
      6'b000000 : _zz_shift_i_0 = shift_i_map_0;
      6'b000001 : _zz_shift_i_0 = shift_i_map_1;
      6'b000010 : _zz_shift_i_0 = shift_i_map_2;
      6'b000011 : _zz_shift_i_0 = shift_i_map_3;
      6'b000100 : _zz_shift_i_0 = shift_i_map_4;
      6'b000101 : _zz_shift_i_0 = shift_i_map_5;
      6'b000110 : _zz_shift_i_0 = shift_i_map_6;
      6'b000111 : _zz_shift_i_0 = shift_i_map_7;
      6'b001000 : _zz_shift_i_0 = shift_i_map_8;
      6'b001001 : _zz_shift_i_0 = shift_i_map_9;
      6'b001010 : _zz_shift_i_0 = shift_i_map_10;
      6'b001011 : _zz_shift_i_0 = shift_i_map_11;
      6'b001100 : _zz_shift_i_0 = shift_i_map_12;
      6'b001101 : _zz_shift_i_0 = shift_i_map_13;
      6'b001110 : _zz_shift_i_0 = shift_i_map_14;
      6'b001111 : _zz_shift_i_0 = shift_i_map_15;
      6'b010000 : _zz_shift_i_0 = shift_i_map_16;
      6'b010001 : _zz_shift_i_0 = shift_i_map_17;
      6'b010010 : _zz_shift_i_0 = shift_i_map_18;
      6'b010011 : _zz_shift_i_0 = shift_i_map_19;
      6'b010100 : _zz_shift_i_0 = shift_i_map_20;
      6'b010101 : _zz_shift_i_0 = shift_i_map_21;
      6'b010110 : _zz_shift_i_0 = shift_i_map_22;
      6'b010111 : _zz_shift_i_0 = shift_i_map_23;
      6'b011000 : _zz_shift_i_0 = shift_i_map_24;
      6'b011001 : _zz_shift_i_0 = shift_i_map_25;
      6'b011010 : _zz_shift_i_0 = shift_i_map_26;
      6'b011011 : _zz_shift_i_0 = shift_i_map_27;
      6'b011100 : _zz_shift_i_0 = shift_i_map_28;
      6'b011101 : _zz_shift_i_0 = shift_i_map_29;
      6'b011110 : _zz_shift_i_0 = shift_i_map_30;
      6'b011111 : _zz_shift_i_0 = shift_i_map_31;
      6'b100000 : _zz_shift_i_0 = shift_i_map_32;
      6'b100001 : _zz_shift_i_0 = shift_i_map_33;
      6'b100010 : _zz_shift_i_0 = shift_i_map_34;
      6'b100011 : _zz_shift_i_0 = shift_i_map_35;
      6'b100100 : _zz_shift_i_0 = shift_i_map_36;
      6'b100101 : _zz_shift_i_0 = shift_i_map_37;
      6'b100110 : _zz_shift_i_0 = shift_i_map_38;
      6'b100111 : _zz_shift_i_0 = shift_i_map_39;
      6'b101000 : _zz_shift_i_0 = shift_i_map_40;
      6'b101001 : _zz_shift_i_0 = shift_i_map_41;
      6'b101010 : _zz_shift_i_0 = shift_i_map_42;
      6'b101011 : _zz_shift_i_0 = shift_i_map_43;
      6'b101100 : _zz_shift_i_0 = shift_i_map_44;
      6'b101101 : _zz_shift_i_0 = shift_i_map_45;
      6'b101110 : _zz_shift_i_0 = shift_i_map_46;
      6'b101111 : _zz_shift_i_0 = shift_i_map_47;
      6'b110000 : _zz_shift_i_0 = shift_i_map_48;
      6'b110001 : _zz_shift_i_0 = shift_i_map_49;
      6'b110010 : _zz_shift_i_0 = shift_i_map_50;
      6'b110011 : _zz_shift_i_0 = shift_i_map_51;
      6'b110100 : _zz_shift_i_0 = shift_i_map_52;
      6'b110101 : _zz_shift_i_0 = shift_i_map_53;
      6'b110110 : _zz_shift_i_0 = shift_i_map_54;
      6'b110111 : _zz_shift_i_0 = shift_i_map_55;
      6'b111000 : _zz_shift_i_0 = shift_i_map_56;
      6'b111001 : _zz_shift_i_0 = shift_i_map_57;
      6'b111010 : _zz_shift_i_0 = shift_i_map_58;
      6'b111011 : _zz_shift_i_0 = shift_i_map_59;
      6'b111100 : _zz_shift_i_0 = shift_i_map_60;
      6'b111101 : _zz_shift_i_0 = shift_i_map_61;
      6'b111110 : _zz_shift_i_0 = shift_i_map_62;
      default : _zz_shift_i_0 = shift_i_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_0_1)
      6'b000000 : _zz_shift_q_0 = shift_q_map_0;
      6'b000001 : _zz_shift_q_0 = shift_q_map_1;
      6'b000010 : _zz_shift_q_0 = shift_q_map_2;
      6'b000011 : _zz_shift_q_0 = shift_q_map_3;
      6'b000100 : _zz_shift_q_0 = shift_q_map_4;
      6'b000101 : _zz_shift_q_0 = shift_q_map_5;
      6'b000110 : _zz_shift_q_0 = shift_q_map_6;
      6'b000111 : _zz_shift_q_0 = shift_q_map_7;
      6'b001000 : _zz_shift_q_0 = shift_q_map_8;
      6'b001001 : _zz_shift_q_0 = shift_q_map_9;
      6'b001010 : _zz_shift_q_0 = shift_q_map_10;
      6'b001011 : _zz_shift_q_0 = shift_q_map_11;
      6'b001100 : _zz_shift_q_0 = shift_q_map_12;
      6'b001101 : _zz_shift_q_0 = shift_q_map_13;
      6'b001110 : _zz_shift_q_0 = shift_q_map_14;
      6'b001111 : _zz_shift_q_0 = shift_q_map_15;
      6'b010000 : _zz_shift_q_0 = shift_q_map_16;
      6'b010001 : _zz_shift_q_0 = shift_q_map_17;
      6'b010010 : _zz_shift_q_0 = shift_q_map_18;
      6'b010011 : _zz_shift_q_0 = shift_q_map_19;
      6'b010100 : _zz_shift_q_0 = shift_q_map_20;
      6'b010101 : _zz_shift_q_0 = shift_q_map_21;
      6'b010110 : _zz_shift_q_0 = shift_q_map_22;
      6'b010111 : _zz_shift_q_0 = shift_q_map_23;
      6'b011000 : _zz_shift_q_0 = shift_q_map_24;
      6'b011001 : _zz_shift_q_0 = shift_q_map_25;
      6'b011010 : _zz_shift_q_0 = shift_q_map_26;
      6'b011011 : _zz_shift_q_0 = shift_q_map_27;
      6'b011100 : _zz_shift_q_0 = shift_q_map_28;
      6'b011101 : _zz_shift_q_0 = shift_q_map_29;
      6'b011110 : _zz_shift_q_0 = shift_q_map_30;
      6'b011111 : _zz_shift_q_0 = shift_q_map_31;
      6'b100000 : _zz_shift_q_0 = shift_q_map_32;
      6'b100001 : _zz_shift_q_0 = shift_q_map_33;
      6'b100010 : _zz_shift_q_0 = shift_q_map_34;
      6'b100011 : _zz_shift_q_0 = shift_q_map_35;
      6'b100100 : _zz_shift_q_0 = shift_q_map_36;
      6'b100101 : _zz_shift_q_0 = shift_q_map_37;
      6'b100110 : _zz_shift_q_0 = shift_q_map_38;
      6'b100111 : _zz_shift_q_0 = shift_q_map_39;
      6'b101000 : _zz_shift_q_0 = shift_q_map_40;
      6'b101001 : _zz_shift_q_0 = shift_q_map_41;
      6'b101010 : _zz_shift_q_0 = shift_q_map_42;
      6'b101011 : _zz_shift_q_0 = shift_q_map_43;
      6'b101100 : _zz_shift_q_0 = shift_q_map_44;
      6'b101101 : _zz_shift_q_0 = shift_q_map_45;
      6'b101110 : _zz_shift_q_0 = shift_q_map_46;
      6'b101111 : _zz_shift_q_0 = shift_q_map_47;
      6'b110000 : _zz_shift_q_0 = shift_q_map_48;
      6'b110001 : _zz_shift_q_0 = shift_q_map_49;
      6'b110010 : _zz_shift_q_0 = shift_q_map_50;
      6'b110011 : _zz_shift_q_0 = shift_q_map_51;
      6'b110100 : _zz_shift_q_0 = shift_q_map_52;
      6'b110101 : _zz_shift_q_0 = shift_q_map_53;
      6'b110110 : _zz_shift_q_0 = shift_q_map_54;
      6'b110111 : _zz_shift_q_0 = shift_q_map_55;
      6'b111000 : _zz_shift_q_0 = shift_q_map_56;
      6'b111001 : _zz_shift_q_0 = shift_q_map_57;
      6'b111010 : _zz_shift_q_0 = shift_q_map_58;
      6'b111011 : _zz_shift_q_0 = shift_q_map_59;
      6'b111100 : _zz_shift_q_0 = shift_q_map_60;
      6'b111101 : _zz_shift_q_0 = shift_q_map_61;
      6'b111110 : _zz_shift_q_0 = shift_q_map_62;
      default : _zz_shift_q_0 = shift_q_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_1_1)
      6'b000000 : _zz_shift_i_1 = shift_i_map_0;
      6'b000001 : _zz_shift_i_1 = shift_i_map_1;
      6'b000010 : _zz_shift_i_1 = shift_i_map_2;
      6'b000011 : _zz_shift_i_1 = shift_i_map_3;
      6'b000100 : _zz_shift_i_1 = shift_i_map_4;
      6'b000101 : _zz_shift_i_1 = shift_i_map_5;
      6'b000110 : _zz_shift_i_1 = shift_i_map_6;
      6'b000111 : _zz_shift_i_1 = shift_i_map_7;
      6'b001000 : _zz_shift_i_1 = shift_i_map_8;
      6'b001001 : _zz_shift_i_1 = shift_i_map_9;
      6'b001010 : _zz_shift_i_1 = shift_i_map_10;
      6'b001011 : _zz_shift_i_1 = shift_i_map_11;
      6'b001100 : _zz_shift_i_1 = shift_i_map_12;
      6'b001101 : _zz_shift_i_1 = shift_i_map_13;
      6'b001110 : _zz_shift_i_1 = shift_i_map_14;
      6'b001111 : _zz_shift_i_1 = shift_i_map_15;
      6'b010000 : _zz_shift_i_1 = shift_i_map_16;
      6'b010001 : _zz_shift_i_1 = shift_i_map_17;
      6'b010010 : _zz_shift_i_1 = shift_i_map_18;
      6'b010011 : _zz_shift_i_1 = shift_i_map_19;
      6'b010100 : _zz_shift_i_1 = shift_i_map_20;
      6'b010101 : _zz_shift_i_1 = shift_i_map_21;
      6'b010110 : _zz_shift_i_1 = shift_i_map_22;
      6'b010111 : _zz_shift_i_1 = shift_i_map_23;
      6'b011000 : _zz_shift_i_1 = shift_i_map_24;
      6'b011001 : _zz_shift_i_1 = shift_i_map_25;
      6'b011010 : _zz_shift_i_1 = shift_i_map_26;
      6'b011011 : _zz_shift_i_1 = shift_i_map_27;
      6'b011100 : _zz_shift_i_1 = shift_i_map_28;
      6'b011101 : _zz_shift_i_1 = shift_i_map_29;
      6'b011110 : _zz_shift_i_1 = shift_i_map_30;
      6'b011111 : _zz_shift_i_1 = shift_i_map_31;
      6'b100000 : _zz_shift_i_1 = shift_i_map_32;
      6'b100001 : _zz_shift_i_1 = shift_i_map_33;
      6'b100010 : _zz_shift_i_1 = shift_i_map_34;
      6'b100011 : _zz_shift_i_1 = shift_i_map_35;
      6'b100100 : _zz_shift_i_1 = shift_i_map_36;
      6'b100101 : _zz_shift_i_1 = shift_i_map_37;
      6'b100110 : _zz_shift_i_1 = shift_i_map_38;
      6'b100111 : _zz_shift_i_1 = shift_i_map_39;
      6'b101000 : _zz_shift_i_1 = shift_i_map_40;
      6'b101001 : _zz_shift_i_1 = shift_i_map_41;
      6'b101010 : _zz_shift_i_1 = shift_i_map_42;
      6'b101011 : _zz_shift_i_1 = shift_i_map_43;
      6'b101100 : _zz_shift_i_1 = shift_i_map_44;
      6'b101101 : _zz_shift_i_1 = shift_i_map_45;
      6'b101110 : _zz_shift_i_1 = shift_i_map_46;
      6'b101111 : _zz_shift_i_1 = shift_i_map_47;
      6'b110000 : _zz_shift_i_1 = shift_i_map_48;
      6'b110001 : _zz_shift_i_1 = shift_i_map_49;
      6'b110010 : _zz_shift_i_1 = shift_i_map_50;
      6'b110011 : _zz_shift_i_1 = shift_i_map_51;
      6'b110100 : _zz_shift_i_1 = shift_i_map_52;
      6'b110101 : _zz_shift_i_1 = shift_i_map_53;
      6'b110110 : _zz_shift_i_1 = shift_i_map_54;
      6'b110111 : _zz_shift_i_1 = shift_i_map_55;
      6'b111000 : _zz_shift_i_1 = shift_i_map_56;
      6'b111001 : _zz_shift_i_1 = shift_i_map_57;
      6'b111010 : _zz_shift_i_1 = shift_i_map_58;
      6'b111011 : _zz_shift_i_1 = shift_i_map_59;
      6'b111100 : _zz_shift_i_1 = shift_i_map_60;
      6'b111101 : _zz_shift_i_1 = shift_i_map_61;
      6'b111110 : _zz_shift_i_1 = shift_i_map_62;
      default : _zz_shift_i_1 = shift_i_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_1_1)
      6'b000000 : _zz_shift_q_1 = shift_q_map_0;
      6'b000001 : _zz_shift_q_1 = shift_q_map_1;
      6'b000010 : _zz_shift_q_1 = shift_q_map_2;
      6'b000011 : _zz_shift_q_1 = shift_q_map_3;
      6'b000100 : _zz_shift_q_1 = shift_q_map_4;
      6'b000101 : _zz_shift_q_1 = shift_q_map_5;
      6'b000110 : _zz_shift_q_1 = shift_q_map_6;
      6'b000111 : _zz_shift_q_1 = shift_q_map_7;
      6'b001000 : _zz_shift_q_1 = shift_q_map_8;
      6'b001001 : _zz_shift_q_1 = shift_q_map_9;
      6'b001010 : _zz_shift_q_1 = shift_q_map_10;
      6'b001011 : _zz_shift_q_1 = shift_q_map_11;
      6'b001100 : _zz_shift_q_1 = shift_q_map_12;
      6'b001101 : _zz_shift_q_1 = shift_q_map_13;
      6'b001110 : _zz_shift_q_1 = shift_q_map_14;
      6'b001111 : _zz_shift_q_1 = shift_q_map_15;
      6'b010000 : _zz_shift_q_1 = shift_q_map_16;
      6'b010001 : _zz_shift_q_1 = shift_q_map_17;
      6'b010010 : _zz_shift_q_1 = shift_q_map_18;
      6'b010011 : _zz_shift_q_1 = shift_q_map_19;
      6'b010100 : _zz_shift_q_1 = shift_q_map_20;
      6'b010101 : _zz_shift_q_1 = shift_q_map_21;
      6'b010110 : _zz_shift_q_1 = shift_q_map_22;
      6'b010111 : _zz_shift_q_1 = shift_q_map_23;
      6'b011000 : _zz_shift_q_1 = shift_q_map_24;
      6'b011001 : _zz_shift_q_1 = shift_q_map_25;
      6'b011010 : _zz_shift_q_1 = shift_q_map_26;
      6'b011011 : _zz_shift_q_1 = shift_q_map_27;
      6'b011100 : _zz_shift_q_1 = shift_q_map_28;
      6'b011101 : _zz_shift_q_1 = shift_q_map_29;
      6'b011110 : _zz_shift_q_1 = shift_q_map_30;
      6'b011111 : _zz_shift_q_1 = shift_q_map_31;
      6'b100000 : _zz_shift_q_1 = shift_q_map_32;
      6'b100001 : _zz_shift_q_1 = shift_q_map_33;
      6'b100010 : _zz_shift_q_1 = shift_q_map_34;
      6'b100011 : _zz_shift_q_1 = shift_q_map_35;
      6'b100100 : _zz_shift_q_1 = shift_q_map_36;
      6'b100101 : _zz_shift_q_1 = shift_q_map_37;
      6'b100110 : _zz_shift_q_1 = shift_q_map_38;
      6'b100111 : _zz_shift_q_1 = shift_q_map_39;
      6'b101000 : _zz_shift_q_1 = shift_q_map_40;
      6'b101001 : _zz_shift_q_1 = shift_q_map_41;
      6'b101010 : _zz_shift_q_1 = shift_q_map_42;
      6'b101011 : _zz_shift_q_1 = shift_q_map_43;
      6'b101100 : _zz_shift_q_1 = shift_q_map_44;
      6'b101101 : _zz_shift_q_1 = shift_q_map_45;
      6'b101110 : _zz_shift_q_1 = shift_q_map_46;
      6'b101111 : _zz_shift_q_1 = shift_q_map_47;
      6'b110000 : _zz_shift_q_1 = shift_q_map_48;
      6'b110001 : _zz_shift_q_1 = shift_q_map_49;
      6'b110010 : _zz_shift_q_1 = shift_q_map_50;
      6'b110011 : _zz_shift_q_1 = shift_q_map_51;
      6'b110100 : _zz_shift_q_1 = shift_q_map_52;
      6'b110101 : _zz_shift_q_1 = shift_q_map_53;
      6'b110110 : _zz_shift_q_1 = shift_q_map_54;
      6'b110111 : _zz_shift_q_1 = shift_q_map_55;
      6'b111000 : _zz_shift_q_1 = shift_q_map_56;
      6'b111001 : _zz_shift_q_1 = shift_q_map_57;
      6'b111010 : _zz_shift_q_1 = shift_q_map_58;
      6'b111011 : _zz_shift_q_1 = shift_q_map_59;
      6'b111100 : _zz_shift_q_1 = shift_q_map_60;
      6'b111101 : _zz_shift_q_1 = shift_q_map_61;
      6'b111110 : _zz_shift_q_1 = shift_q_map_62;
      default : _zz_shift_q_1 = shift_q_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_2_1)
      6'b000000 : _zz_shift_i_2 = shift_i_map_0;
      6'b000001 : _zz_shift_i_2 = shift_i_map_1;
      6'b000010 : _zz_shift_i_2 = shift_i_map_2;
      6'b000011 : _zz_shift_i_2 = shift_i_map_3;
      6'b000100 : _zz_shift_i_2 = shift_i_map_4;
      6'b000101 : _zz_shift_i_2 = shift_i_map_5;
      6'b000110 : _zz_shift_i_2 = shift_i_map_6;
      6'b000111 : _zz_shift_i_2 = shift_i_map_7;
      6'b001000 : _zz_shift_i_2 = shift_i_map_8;
      6'b001001 : _zz_shift_i_2 = shift_i_map_9;
      6'b001010 : _zz_shift_i_2 = shift_i_map_10;
      6'b001011 : _zz_shift_i_2 = shift_i_map_11;
      6'b001100 : _zz_shift_i_2 = shift_i_map_12;
      6'b001101 : _zz_shift_i_2 = shift_i_map_13;
      6'b001110 : _zz_shift_i_2 = shift_i_map_14;
      6'b001111 : _zz_shift_i_2 = shift_i_map_15;
      6'b010000 : _zz_shift_i_2 = shift_i_map_16;
      6'b010001 : _zz_shift_i_2 = shift_i_map_17;
      6'b010010 : _zz_shift_i_2 = shift_i_map_18;
      6'b010011 : _zz_shift_i_2 = shift_i_map_19;
      6'b010100 : _zz_shift_i_2 = shift_i_map_20;
      6'b010101 : _zz_shift_i_2 = shift_i_map_21;
      6'b010110 : _zz_shift_i_2 = shift_i_map_22;
      6'b010111 : _zz_shift_i_2 = shift_i_map_23;
      6'b011000 : _zz_shift_i_2 = shift_i_map_24;
      6'b011001 : _zz_shift_i_2 = shift_i_map_25;
      6'b011010 : _zz_shift_i_2 = shift_i_map_26;
      6'b011011 : _zz_shift_i_2 = shift_i_map_27;
      6'b011100 : _zz_shift_i_2 = shift_i_map_28;
      6'b011101 : _zz_shift_i_2 = shift_i_map_29;
      6'b011110 : _zz_shift_i_2 = shift_i_map_30;
      6'b011111 : _zz_shift_i_2 = shift_i_map_31;
      6'b100000 : _zz_shift_i_2 = shift_i_map_32;
      6'b100001 : _zz_shift_i_2 = shift_i_map_33;
      6'b100010 : _zz_shift_i_2 = shift_i_map_34;
      6'b100011 : _zz_shift_i_2 = shift_i_map_35;
      6'b100100 : _zz_shift_i_2 = shift_i_map_36;
      6'b100101 : _zz_shift_i_2 = shift_i_map_37;
      6'b100110 : _zz_shift_i_2 = shift_i_map_38;
      6'b100111 : _zz_shift_i_2 = shift_i_map_39;
      6'b101000 : _zz_shift_i_2 = shift_i_map_40;
      6'b101001 : _zz_shift_i_2 = shift_i_map_41;
      6'b101010 : _zz_shift_i_2 = shift_i_map_42;
      6'b101011 : _zz_shift_i_2 = shift_i_map_43;
      6'b101100 : _zz_shift_i_2 = shift_i_map_44;
      6'b101101 : _zz_shift_i_2 = shift_i_map_45;
      6'b101110 : _zz_shift_i_2 = shift_i_map_46;
      6'b101111 : _zz_shift_i_2 = shift_i_map_47;
      6'b110000 : _zz_shift_i_2 = shift_i_map_48;
      6'b110001 : _zz_shift_i_2 = shift_i_map_49;
      6'b110010 : _zz_shift_i_2 = shift_i_map_50;
      6'b110011 : _zz_shift_i_2 = shift_i_map_51;
      6'b110100 : _zz_shift_i_2 = shift_i_map_52;
      6'b110101 : _zz_shift_i_2 = shift_i_map_53;
      6'b110110 : _zz_shift_i_2 = shift_i_map_54;
      6'b110111 : _zz_shift_i_2 = shift_i_map_55;
      6'b111000 : _zz_shift_i_2 = shift_i_map_56;
      6'b111001 : _zz_shift_i_2 = shift_i_map_57;
      6'b111010 : _zz_shift_i_2 = shift_i_map_58;
      6'b111011 : _zz_shift_i_2 = shift_i_map_59;
      6'b111100 : _zz_shift_i_2 = shift_i_map_60;
      6'b111101 : _zz_shift_i_2 = shift_i_map_61;
      6'b111110 : _zz_shift_i_2 = shift_i_map_62;
      default : _zz_shift_i_2 = shift_i_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_2_1)
      6'b000000 : _zz_shift_q_2 = shift_q_map_0;
      6'b000001 : _zz_shift_q_2 = shift_q_map_1;
      6'b000010 : _zz_shift_q_2 = shift_q_map_2;
      6'b000011 : _zz_shift_q_2 = shift_q_map_3;
      6'b000100 : _zz_shift_q_2 = shift_q_map_4;
      6'b000101 : _zz_shift_q_2 = shift_q_map_5;
      6'b000110 : _zz_shift_q_2 = shift_q_map_6;
      6'b000111 : _zz_shift_q_2 = shift_q_map_7;
      6'b001000 : _zz_shift_q_2 = shift_q_map_8;
      6'b001001 : _zz_shift_q_2 = shift_q_map_9;
      6'b001010 : _zz_shift_q_2 = shift_q_map_10;
      6'b001011 : _zz_shift_q_2 = shift_q_map_11;
      6'b001100 : _zz_shift_q_2 = shift_q_map_12;
      6'b001101 : _zz_shift_q_2 = shift_q_map_13;
      6'b001110 : _zz_shift_q_2 = shift_q_map_14;
      6'b001111 : _zz_shift_q_2 = shift_q_map_15;
      6'b010000 : _zz_shift_q_2 = shift_q_map_16;
      6'b010001 : _zz_shift_q_2 = shift_q_map_17;
      6'b010010 : _zz_shift_q_2 = shift_q_map_18;
      6'b010011 : _zz_shift_q_2 = shift_q_map_19;
      6'b010100 : _zz_shift_q_2 = shift_q_map_20;
      6'b010101 : _zz_shift_q_2 = shift_q_map_21;
      6'b010110 : _zz_shift_q_2 = shift_q_map_22;
      6'b010111 : _zz_shift_q_2 = shift_q_map_23;
      6'b011000 : _zz_shift_q_2 = shift_q_map_24;
      6'b011001 : _zz_shift_q_2 = shift_q_map_25;
      6'b011010 : _zz_shift_q_2 = shift_q_map_26;
      6'b011011 : _zz_shift_q_2 = shift_q_map_27;
      6'b011100 : _zz_shift_q_2 = shift_q_map_28;
      6'b011101 : _zz_shift_q_2 = shift_q_map_29;
      6'b011110 : _zz_shift_q_2 = shift_q_map_30;
      6'b011111 : _zz_shift_q_2 = shift_q_map_31;
      6'b100000 : _zz_shift_q_2 = shift_q_map_32;
      6'b100001 : _zz_shift_q_2 = shift_q_map_33;
      6'b100010 : _zz_shift_q_2 = shift_q_map_34;
      6'b100011 : _zz_shift_q_2 = shift_q_map_35;
      6'b100100 : _zz_shift_q_2 = shift_q_map_36;
      6'b100101 : _zz_shift_q_2 = shift_q_map_37;
      6'b100110 : _zz_shift_q_2 = shift_q_map_38;
      6'b100111 : _zz_shift_q_2 = shift_q_map_39;
      6'b101000 : _zz_shift_q_2 = shift_q_map_40;
      6'b101001 : _zz_shift_q_2 = shift_q_map_41;
      6'b101010 : _zz_shift_q_2 = shift_q_map_42;
      6'b101011 : _zz_shift_q_2 = shift_q_map_43;
      6'b101100 : _zz_shift_q_2 = shift_q_map_44;
      6'b101101 : _zz_shift_q_2 = shift_q_map_45;
      6'b101110 : _zz_shift_q_2 = shift_q_map_46;
      6'b101111 : _zz_shift_q_2 = shift_q_map_47;
      6'b110000 : _zz_shift_q_2 = shift_q_map_48;
      6'b110001 : _zz_shift_q_2 = shift_q_map_49;
      6'b110010 : _zz_shift_q_2 = shift_q_map_50;
      6'b110011 : _zz_shift_q_2 = shift_q_map_51;
      6'b110100 : _zz_shift_q_2 = shift_q_map_52;
      6'b110101 : _zz_shift_q_2 = shift_q_map_53;
      6'b110110 : _zz_shift_q_2 = shift_q_map_54;
      6'b110111 : _zz_shift_q_2 = shift_q_map_55;
      6'b111000 : _zz_shift_q_2 = shift_q_map_56;
      6'b111001 : _zz_shift_q_2 = shift_q_map_57;
      6'b111010 : _zz_shift_q_2 = shift_q_map_58;
      6'b111011 : _zz_shift_q_2 = shift_q_map_59;
      6'b111100 : _zz_shift_q_2 = shift_q_map_60;
      6'b111101 : _zz_shift_q_2 = shift_q_map_61;
      6'b111110 : _zz_shift_q_2 = shift_q_map_62;
      default : _zz_shift_q_2 = shift_q_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_3_1)
      6'b000000 : _zz_shift_i_3 = shift_i_map_0;
      6'b000001 : _zz_shift_i_3 = shift_i_map_1;
      6'b000010 : _zz_shift_i_3 = shift_i_map_2;
      6'b000011 : _zz_shift_i_3 = shift_i_map_3;
      6'b000100 : _zz_shift_i_3 = shift_i_map_4;
      6'b000101 : _zz_shift_i_3 = shift_i_map_5;
      6'b000110 : _zz_shift_i_3 = shift_i_map_6;
      6'b000111 : _zz_shift_i_3 = shift_i_map_7;
      6'b001000 : _zz_shift_i_3 = shift_i_map_8;
      6'b001001 : _zz_shift_i_3 = shift_i_map_9;
      6'b001010 : _zz_shift_i_3 = shift_i_map_10;
      6'b001011 : _zz_shift_i_3 = shift_i_map_11;
      6'b001100 : _zz_shift_i_3 = shift_i_map_12;
      6'b001101 : _zz_shift_i_3 = shift_i_map_13;
      6'b001110 : _zz_shift_i_3 = shift_i_map_14;
      6'b001111 : _zz_shift_i_3 = shift_i_map_15;
      6'b010000 : _zz_shift_i_3 = shift_i_map_16;
      6'b010001 : _zz_shift_i_3 = shift_i_map_17;
      6'b010010 : _zz_shift_i_3 = shift_i_map_18;
      6'b010011 : _zz_shift_i_3 = shift_i_map_19;
      6'b010100 : _zz_shift_i_3 = shift_i_map_20;
      6'b010101 : _zz_shift_i_3 = shift_i_map_21;
      6'b010110 : _zz_shift_i_3 = shift_i_map_22;
      6'b010111 : _zz_shift_i_3 = shift_i_map_23;
      6'b011000 : _zz_shift_i_3 = shift_i_map_24;
      6'b011001 : _zz_shift_i_3 = shift_i_map_25;
      6'b011010 : _zz_shift_i_3 = shift_i_map_26;
      6'b011011 : _zz_shift_i_3 = shift_i_map_27;
      6'b011100 : _zz_shift_i_3 = shift_i_map_28;
      6'b011101 : _zz_shift_i_3 = shift_i_map_29;
      6'b011110 : _zz_shift_i_3 = shift_i_map_30;
      6'b011111 : _zz_shift_i_3 = shift_i_map_31;
      6'b100000 : _zz_shift_i_3 = shift_i_map_32;
      6'b100001 : _zz_shift_i_3 = shift_i_map_33;
      6'b100010 : _zz_shift_i_3 = shift_i_map_34;
      6'b100011 : _zz_shift_i_3 = shift_i_map_35;
      6'b100100 : _zz_shift_i_3 = shift_i_map_36;
      6'b100101 : _zz_shift_i_3 = shift_i_map_37;
      6'b100110 : _zz_shift_i_3 = shift_i_map_38;
      6'b100111 : _zz_shift_i_3 = shift_i_map_39;
      6'b101000 : _zz_shift_i_3 = shift_i_map_40;
      6'b101001 : _zz_shift_i_3 = shift_i_map_41;
      6'b101010 : _zz_shift_i_3 = shift_i_map_42;
      6'b101011 : _zz_shift_i_3 = shift_i_map_43;
      6'b101100 : _zz_shift_i_3 = shift_i_map_44;
      6'b101101 : _zz_shift_i_3 = shift_i_map_45;
      6'b101110 : _zz_shift_i_3 = shift_i_map_46;
      6'b101111 : _zz_shift_i_3 = shift_i_map_47;
      6'b110000 : _zz_shift_i_3 = shift_i_map_48;
      6'b110001 : _zz_shift_i_3 = shift_i_map_49;
      6'b110010 : _zz_shift_i_3 = shift_i_map_50;
      6'b110011 : _zz_shift_i_3 = shift_i_map_51;
      6'b110100 : _zz_shift_i_3 = shift_i_map_52;
      6'b110101 : _zz_shift_i_3 = shift_i_map_53;
      6'b110110 : _zz_shift_i_3 = shift_i_map_54;
      6'b110111 : _zz_shift_i_3 = shift_i_map_55;
      6'b111000 : _zz_shift_i_3 = shift_i_map_56;
      6'b111001 : _zz_shift_i_3 = shift_i_map_57;
      6'b111010 : _zz_shift_i_3 = shift_i_map_58;
      6'b111011 : _zz_shift_i_3 = shift_i_map_59;
      6'b111100 : _zz_shift_i_3 = shift_i_map_60;
      6'b111101 : _zz_shift_i_3 = shift_i_map_61;
      6'b111110 : _zz_shift_i_3 = shift_i_map_62;
      default : _zz_shift_i_3 = shift_i_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_3_1)
      6'b000000 : _zz_shift_q_3 = shift_q_map_0;
      6'b000001 : _zz_shift_q_3 = shift_q_map_1;
      6'b000010 : _zz_shift_q_3 = shift_q_map_2;
      6'b000011 : _zz_shift_q_3 = shift_q_map_3;
      6'b000100 : _zz_shift_q_3 = shift_q_map_4;
      6'b000101 : _zz_shift_q_3 = shift_q_map_5;
      6'b000110 : _zz_shift_q_3 = shift_q_map_6;
      6'b000111 : _zz_shift_q_3 = shift_q_map_7;
      6'b001000 : _zz_shift_q_3 = shift_q_map_8;
      6'b001001 : _zz_shift_q_3 = shift_q_map_9;
      6'b001010 : _zz_shift_q_3 = shift_q_map_10;
      6'b001011 : _zz_shift_q_3 = shift_q_map_11;
      6'b001100 : _zz_shift_q_3 = shift_q_map_12;
      6'b001101 : _zz_shift_q_3 = shift_q_map_13;
      6'b001110 : _zz_shift_q_3 = shift_q_map_14;
      6'b001111 : _zz_shift_q_3 = shift_q_map_15;
      6'b010000 : _zz_shift_q_3 = shift_q_map_16;
      6'b010001 : _zz_shift_q_3 = shift_q_map_17;
      6'b010010 : _zz_shift_q_3 = shift_q_map_18;
      6'b010011 : _zz_shift_q_3 = shift_q_map_19;
      6'b010100 : _zz_shift_q_3 = shift_q_map_20;
      6'b010101 : _zz_shift_q_3 = shift_q_map_21;
      6'b010110 : _zz_shift_q_3 = shift_q_map_22;
      6'b010111 : _zz_shift_q_3 = shift_q_map_23;
      6'b011000 : _zz_shift_q_3 = shift_q_map_24;
      6'b011001 : _zz_shift_q_3 = shift_q_map_25;
      6'b011010 : _zz_shift_q_3 = shift_q_map_26;
      6'b011011 : _zz_shift_q_3 = shift_q_map_27;
      6'b011100 : _zz_shift_q_3 = shift_q_map_28;
      6'b011101 : _zz_shift_q_3 = shift_q_map_29;
      6'b011110 : _zz_shift_q_3 = shift_q_map_30;
      6'b011111 : _zz_shift_q_3 = shift_q_map_31;
      6'b100000 : _zz_shift_q_3 = shift_q_map_32;
      6'b100001 : _zz_shift_q_3 = shift_q_map_33;
      6'b100010 : _zz_shift_q_3 = shift_q_map_34;
      6'b100011 : _zz_shift_q_3 = shift_q_map_35;
      6'b100100 : _zz_shift_q_3 = shift_q_map_36;
      6'b100101 : _zz_shift_q_3 = shift_q_map_37;
      6'b100110 : _zz_shift_q_3 = shift_q_map_38;
      6'b100111 : _zz_shift_q_3 = shift_q_map_39;
      6'b101000 : _zz_shift_q_3 = shift_q_map_40;
      6'b101001 : _zz_shift_q_3 = shift_q_map_41;
      6'b101010 : _zz_shift_q_3 = shift_q_map_42;
      6'b101011 : _zz_shift_q_3 = shift_q_map_43;
      6'b101100 : _zz_shift_q_3 = shift_q_map_44;
      6'b101101 : _zz_shift_q_3 = shift_q_map_45;
      6'b101110 : _zz_shift_q_3 = shift_q_map_46;
      6'b101111 : _zz_shift_q_3 = shift_q_map_47;
      6'b110000 : _zz_shift_q_3 = shift_q_map_48;
      6'b110001 : _zz_shift_q_3 = shift_q_map_49;
      6'b110010 : _zz_shift_q_3 = shift_q_map_50;
      6'b110011 : _zz_shift_q_3 = shift_q_map_51;
      6'b110100 : _zz_shift_q_3 = shift_q_map_52;
      6'b110101 : _zz_shift_q_3 = shift_q_map_53;
      6'b110110 : _zz_shift_q_3 = shift_q_map_54;
      6'b110111 : _zz_shift_q_3 = shift_q_map_55;
      6'b111000 : _zz_shift_q_3 = shift_q_map_56;
      6'b111001 : _zz_shift_q_3 = shift_q_map_57;
      6'b111010 : _zz_shift_q_3 = shift_q_map_58;
      6'b111011 : _zz_shift_q_3 = shift_q_map_59;
      6'b111100 : _zz_shift_q_3 = shift_q_map_60;
      6'b111101 : _zz_shift_q_3 = shift_q_map_61;
      6'b111110 : _zz_shift_q_3 = shift_q_map_62;
      default : _zz_shift_q_3 = shift_q_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_4_1)
      6'b000000 : _zz_shift_i_4 = shift_i_map_0;
      6'b000001 : _zz_shift_i_4 = shift_i_map_1;
      6'b000010 : _zz_shift_i_4 = shift_i_map_2;
      6'b000011 : _zz_shift_i_4 = shift_i_map_3;
      6'b000100 : _zz_shift_i_4 = shift_i_map_4;
      6'b000101 : _zz_shift_i_4 = shift_i_map_5;
      6'b000110 : _zz_shift_i_4 = shift_i_map_6;
      6'b000111 : _zz_shift_i_4 = shift_i_map_7;
      6'b001000 : _zz_shift_i_4 = shift_i_map_8;
      6'b001001 : _zz_shift_i_4 = shift_i_map_9;
      6'b001010 : _zz_shift_i_4 = shift_i_map_10;
      6'b001011 : _zz_shift_i_4 = shift_i_map_11;
      6'b001100 : _zz_shift_i_4 = shift_i_map_12;
      6'b001101 : _zz_shift_i_4 = shift_i_map_13;
      6'b001110 : _zz_shift_i_4 = shift_i_map_14;
      6'b001111 : _zz_shift_i_4 = shift_i_map_15;
      6'b010000 : _zz_shift_i_4 = shift_i_map_16;
      6'b010001 : _zz_shift_i_4 = shift_i_map_17;
      6'b010010 : _zz_shift_i_4 = shift_i_map_18;
      6'b010011 : _zz_shift_i_4 = shift_i_map_19;
      6'b010100 : _zz_shift_i_4 = shift_i_map_20;
      6'b010101 : _zz_shift_i_4 = shift_i_map_21;
      6'b010110 : _zz_shift_i_4 = shift_i_map_22;
      6'b010111 : _zz_shift_i_4 = shift_i_map_23;
      6'b011000 : _zz_shift_i_4 = shift_i_map_24;
      6'b011001 : _zz_shift_i_4 = shift_i_map_25;
      6'b011010 : _zz_shift_i_4 = shift_i_map_26;
      6'b011011 : _zz_shift_i_4 = shift_i_map_27;
      6'b011100 : _zz_shift_i_4 = shift_i_map_28;
      6'b011101 : _zz_shift_i_4 = shift_i_map_29;
      6'b011110 : _zz_shift_i_4 = shift_i_map_30;
      6'b011111 : _zz_shift_i_4 = shift_i_map_31;
      6'b100000 : _zz_shift_i_4 = shift_i_map_32;
      6'b100001 : _zz_shift_i_4 = shift_i_map_33;
      6'b100010 : _zz_shift_i_4 = shift_i_map_34;
      6'b100011 : _zz_shift_i_4 = shift_i_map_35;
      6'b100100 : _zz_shift_i_4 = shift_i_map_36;
      6'b100101 : _zz_shift_i_4 = shift_i_map_37;
      6'b100110 : _zz_shift_i_4 = shift_i_map_38;
      6'b100111 : _zz_shift_i_4 = shift_i_map_39;
      6'b101000 : _zz_shift_i_4 = shift_i_map_40;
      6'b101001 : _zz_shift_i_4 = shift_i_map_41;
      6'b101010 : _zz_shift_i_4 = shift_i_map_42;
      6'b101011 : _zz_shift_i_4 = shift_i_map_43;
      6'b101100 : _zz_shift_i_4 = shift_i_map_44;
      6'b101101 : _zz_shift_i_4 = shift_i_map_45;
      6'b101110 : _zz_shift_i_4 = shift_i_map_46;
      6'b101111 : _zz_shift_i_4 = shift_i_map_47;
      6'b110000 : _zz_shift_i_4 = shift_i_map_48;
      6'b110001 : _zz_shift_i_4 = shift_i_map_49;
      6'b110010 : _zz_shift_i_4 = shift_i_map_50;
      6'b110011 : _zz_shift_i_4 = shift_i_map_51;
      6'b110100 : _zz_shift_i_4 = shift_i_map_52;
      6'b110101 : _zz_shift_i_4 = shift_i_map_53;
      6'b110110 : _zz_shift_i_4 = shift_i_map_54;
      6'b110111 : _zz_shift_i_4 = shift_i_map_55;
      6'b111000 : _zz_shift_i_4 = shift_i_map_56;
      6'b111001 : _zz_shift_i_4 = shift_i_map_57;
      6'b111010 : _zz_shift_i_4 = shift_i_map_58;
      6'b111011 : _zz_shift_i_4 = shift_i_map_59;
      6'b111100 : _zz_shift_i_4 = shift_i_map_60;
      6'b111101 : _zz_shift_i_4 = shift_i_map_61;
      6'b111110 : _zz_shift_i_4 = shift_i_map_62;
      default : _zz_shift_i_4 = shift_i_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_4_1)
      6'b000000 : _zz_shift_q_4 = shift_q_map_0;
      6'b000001 : _zz_shift_q_4 = shift_q_map_1;
      6'b000010 : _zz_shift_q_4 = shift_q_map_2;
      6'b000011 : _zz_shift_q_4 = shift_q_map_3;
      6'b000100 : _zz_shift_q_4 = shift_q_map_4;
      6'b000101 : _zz_shift_q_4 = shift_q_map_5;
      6'b000110 : _zz_shift_q_4 = shift_q_map_6;
      6'b000111 : _zz_shift_q_4 = shift_q_map_7;
      6'b001000 : _zz_shift_q_4 = shift_q_map_8;
      6'b001001 : _zz_shift_q_4 = shift_q_map_9;
      6'b001010 : _zz_shift_q_4 = shift_q_map_10;
      6'b001011 : _zz_shift_q_4 = shift_q_map_11;
      6'b001100 : _zz_shift_q_4 = shift_q_map_12;
      6'b001101 : _zz_shift_q_4 = shift_q_map_13;
      6'b001110 : _zz_shift_q_4 = shift_q_map_14;
      6'b001111 : _zz_shift_q_4 = shift_q_map_15;
      6'b010000 : _zz_shift_q_4 = shift_q_map_16;
      6'b010001 : _zz_shift_q_4 = shift_q_map_17;
      6'b010010 : _zz_shift_q_4 = shift_q_map_18;
      6'b010011 : _zz_shift_q_4 = shift_q_map_19;
      6'b010100 : _zz_shift_q_4 = shift_q_map_20;
      6'b010101 : _zz_shift_q_4 = shift_q_map_21;
      6'b010110 : _zz_shift_q_4 = shift_q_map_22;
      6'b010111 : _zz_shift_q_4 = shift_q_map_23;
      6'b011000 : _zz_shift_q_4 = shift_q_map_24;
      6'b011001 : _zz_shift_q_4 = shift_q_map_25;
      6'b011010 : _zz_shift_q_4 = shift_q_map_26;
      6'b011011 : _zz_shift_q_4 = shift_q_map_27;
      6'b011100 : _zz_shift_q_4 = shift_q_map_28;
      6'b011101 : _zz_shift_q_4 = shift_q_map_29;
      6'b011110 : _zz_shift_q_4 = shift_q_map_30;
      6'b011111 : _zz_shift_q_4 = shift_q_map_31;
      6'b100000 : _zz_shift_q_4 = shift_q_map_32;
      6'b100001 : _zz_shift_q_4 = shift_q_map_33;
      6'b100010 : _zz_shift_q_4 = shift_q_map_34;
      6'b100011 : _zz_shift_q_4 = shift_q_map_35;
      6'b100100 : _zz_shift_q_4 = shift_q_map_36;
      6'b100101 : _zz_shift_q_4 = shift_q_map_37;
      6'b100110 : _zz_shift_q_4 = shift_q_map_38;
      6'b100111 : _zz_shift_q_4 = shift_q_map_39;
      6'b101000 : _zz_shift_q_4 = shift_q_map_40;
      6'b101001 : _zz_shift_q_4 = shift_q_map_41;
      6'b101010 : _zz_shift_q_4 = shift_q_map_42;
      6'b101011 : _zz_shift_q_4 = shift_q_map_43;
      6'b101100 : _zz_shift_q_4 = shift_q_map_44;
      6'b101101 : _zz_shift_q_4 = shift_q_map_45;
      6'b101110 : _zz_shift_q_4 = shift_q_map_46;
      6'b101111 : _zz_shift_q_4 = shift_q_map_47;
      6'b110000 : _zz_shift_q_4 = shift_q_map_48;
      6'b110001 : _zz_shift_q_4 = shift_q_map_49;
      6'b110010 : _zz_shift_q_4 = shift_q_map_50;
      6'b110011 : _zz_shift_q_4 = shift_q_map_51;
      6'b110100 : _zz_shift_q_4 = shift_q_map_52;
      6'b110101 : _zz_shift_q_4 = shift_q_map_53;
      6'b110110 : _zz_shift_q_4 = shift_q_map_54;
      6'b110111 : _zz_shift_q_4 = shift_q_map_55;
      6'b111000 : _zz_shift_q_4 = shift_q_map_56;
      6'b111001 : _zz_shift_q_4 = shift_q_map_57;
      6'b111010 : _zz_shift_q_4 = shift_q_map_58;
      6'b111011 : _zz_shift_q_4 = shift_q_map_59;
      6'b111100 : _zz_shift_q_4 = shift_q_map_60;
      6'b111101 : _zz_shift_q_4 = shift_q_map_61;
      6'b111110 : _zz_shift_q_4 = shift_q_map_62;
      default : _zz_shift_q_4 = shift_q_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_5_1)
      6'b000000 : _zz_shift_i_5 = shift_i_map_0;
      6'b000001 : _zz_shift_i_5 = shift_i_map_1;
      6'b000010 : _zz_shift_i_5 = shift_i_map_2;
      6'b000011 : _zz_shift_i_5 = shift_i_map_3;
      6'b000100 : _zz_shift_i_5 = shift_i_map_4;
      6'b000101 : _zz_shift_i_5 = shift_i_map_5;
      6'b000110 : _zz_shift_i_5 = shift_i_map_6;
      6'b000111 : _zz_shift_i_5 = shift_i_map_7;
      6'b001000 : _zz_shift_i_5 = shift_i_map_8;
      6'b001001 : _zz_shift_i_5 = shift_i_map_9;
      6'b001010 : _zz_shift_i_5 = shift_i_map_10;
      6'b001011 : _zz_shift_i_5 = shift_i_map_11;
      6'b001100 : _zz_shift_i_5 = shift_i_map_12;
      6'b001101 : _zz_shift_i_5 = shift_i_map_13;
      6'b001110 : _zz_shift_i_5 = shift_i_map_14;
      6'b001111 : _zz_shift_i_5 = shift_i_map_15;
      6'b010000 : _zz_shift_i_5 = shift_i_map_16;
      6'b010001 : _zz_shift_i_5 = shift_i_map_17;
      6'b010010 : _zz_shift_i_5 = shift_i_map_18;
      6'b010011 : _zz_shift_i_5 = shift_i_map_19;
      6'b010100 : _zz_shift_i_5 = shift_i_map_20;
      6'b010101 : _zz_shift_i_5 = shift_i_map_21;
      6'b010110 : _zz_shift_i_5 = shift_i_map_22;
      6'b010111 : _zz_shift_i_5 = shift_i_map_23;
      6'b011000 : _zz_shift_i_5 = shift_i_map_24;
      6'b011001 : _zz_shift_i_5 = shift_i_map_25;
      6'b011010 : _zz_shift_i_5 = shift_i_map_26;
      6'b011011 : _zz_shift_i_5 = shift_i_map_27;
      6'b011100 : _zz_shift_i_5 = shift_i_map_28;
      6'b011101 : _zz_shift_i_5 = shift_i_map_29;
      6'b011110 : _zz_shift_i_5 = shift_i_map_30;
      6'b011111 : _zz_shift_i_5 = shift_i_map_31;
      6'b100000 : _zz_shift_i_5 = shift_i_map_32;
      6'b100001 : _zz_shift_i_5 = shift_i_map_33;
      6'b100010 : _zz_shift_i_5 = shift_i_map_34;
      6'b100011 : _zz_shift_i_5 = shift_i_map_35;
      6'b100100 : _zz_shift_i_5 = shift_i_map_36;
      6'b100101 : _zz_shift_i_5 = shift_i_map_37;
      6'b100110 : _zz_shift_i_5 = shift_i_map_38;
      6'b100111 : _zz_shift_i_5 = shift_i_map_39;
      6'b101000 : _zz_shift_i_5 = shift_i_map_40;
      6'b101001 : _zz_shift_i_5 = shift_i_map_41;
      6'b101010 : _zz_shift_i_5 = shift_i_map_42;
      6'b101011 : _zz_shift_i_5 = shift_i_map_43;
      6'b101100 : _zz_shift_i_5 = shift_i_map_44;
      6'b101101 : _zz_shift_i_5 = shift_i_map_45;
      6'b101110 : _zz_shift_i_5 = shift_i_map_46;
      6'b101111 : _zz_shift_i_5 = shift_i_map_47;
      6'b110000 : _zz_shift_i_5 = shift_i_map_48;
      6'b110001 : _zz_shift_i_5 = shift_i_map_49;
      6'b110010 : _zz_shift_i_5 = shift_i_map_50;
      6'b110011 : _zz_shift_i_5 = shift_i_map_51;
      6'b110100 : _zz_shift_i_5 = shift_i_map_52;
      6'b110101 : _zz_shift_i_5 = shift_i_map_53;
      6'b110110 : _zz_shift_i_5 = shift_i_map_54;
      6'b110111 : _zz_shift_i_5 = shift_i_map_55;
      6'b111000 : _zz_shift_i_5 = shift_i_map_56;
      6'b111001 : _zz_shift_i_5 = shift_i_map_57;
      6'b111010 : _zz_shift_i_5 = shift_i_map_58;
      6'b111011 : _zz_shift_i_5 = shift_i_map_59;
      6'b111100 : _zz_shift_i_5 = shift_i_map_60;
      6'b111101 : _zz_shift_i_5 = shift_i_map_61;
      6'b111110 : _zz_shift_i_5 = shift_i_map_62;
      default : _zz_shift_i_5 = shift_i_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_5_1)
      6'b000000 : _zz_shift_q_5 = shift_q_map_0;
      6'b000001 : _zz_shift_q_5 = shift_q_map_1;
      6'b000010 : _zz_shift_q_5 = shift_q_map_2;
      6'b000011 : _zz_shift_q_5 = shift_q_map_3;
      6'b000100 : _zz_shift_q_5 = shift_q_map_4;
      6'b000101 : _zz_shift_q_5 = shift_q_map_5;
      6'b000110 : _zz_shift_q_5 = shift_q_map_6;
      6'b000111 : _zz_shift_q_5 = shift_q_map_7;
      6'b001000 : _zz_shift_q_5 = shift_q_map_8;
      6'b001001 : _zz_shift_q_5 = shift_q_map_9;
      6'b001010 : _zz_shift_q_5 = shift_q_map_10;
      6'b001011 : _zz_shift_q_5 = shift_q_map_11;
      6'b001100 : _zz_shift_q_5 = shift_q_map_12;
      6'b001101 : _zz_shift_q_5 = shift_q_map_13;
      6'b001110 : _zz_shift_q_5 = shift_q_map_14;
      6'b001111 : _zz_shift_q_5 = shift_q_map_15;
      6'b010000 : _zz_shift_q_5 = shift_q_map_16;
      6'b010001 : _zz_shift_q_5 = shift_q_map_17;
      6'b010010 : _zz_shift_q_5 = shift_q_map_18;
      6'b010011 : _zz_shift_q_5 = shift_q_map_19;
      6'b010100 : _zz_shift_q_5 = shift_q_map_20;
      6'b010101 : _zz_shift_q_5 = shift_q_map_21;
      6'b010110 : _zz_shift_q_5 = shift_q_map_22;
      6'b010111 : _zz_shift_q_5 = shift_q_map_23;
      6'b011000 : _zz_shift_q_5 = shift_q_map_24;
      6'b011001 : _zz_shift_q_5 = shift_q_map_25;
      6'b011010 : _zz_shift_q_5 = shift_q_map_26;
      6'b011011 : _zz_shift_q_5 = shift_q_map_27;
      6'b011100 : _zz_shift_q_5 = shift_q_map_28;
      6'b011101 : _zz_shift_q_5 = shift_q_map_29;
      6'b011110 : _zz_shift_q_5 = shift_q_map_30;
      6'b011111 : _zz_shift_q_5 = shift_q_map_31;
      6'b100000 : _zz_shift_q_5 = shift_q_map_32;
      6'b100001 : _zz_shift_q_5 = shift_q_map_33;
      6'b100010 : _zz_shift_q_5 = shift_q_map_34;
      6'b100011 : _zz_shift_q_5 = shift_q_map_35;
      6'b100100 : _zz_shift_q_5 = shift_q_map_36;
      6'b100101 : _zz_shift_q_5 = shift_q_map_37;
      6'b100110 : _zz_shift_q_5 = shift_q_map_38;
      6'b100111 : _zz_shift_q_5 = shift_q_map_39;
      6'b101000 : _zz_shift_q_5 = shift_q_map_40;
      6'b101001 : _zz_shift_q_5 = shift_q_map_41;
      6'b101010 : _zz_shift_q_5 = shift_q_map_42;
      6'b101011 : _zz_shift_q_5 = shift_q_map_43;
      6'b101100 : _zz_shift_q_5 = shift_q_map_44;
      6'b101101 : _zz_shift_q_5 = shift_q_map_45;
      6'b101110 : _zz_shift_q_5 = shift_q_map_46;
      6'b101111 : _zz_shift_q_5 = shift_q_map_47;
      6'b110000 : _zz_shift_q_5 = shift_q_map_48;
      6'b110001 : _zz_shift_q_5 = shift_q_map_49;
      6'b110010 : _zz_shift_q_5 = shift_q_map_50;
      6'b110011 : _zz_shift_q_5 = shift_q_map_51;
      6'b110100 : _zz_shift_q_5 = shift_q_map_52;
      6'b110101 : _zz_shift_q_5 = shift_q_map_53;
      6'b110110 : _zz_shift_q_5 = shift_q_map_54;
      6'b110111 : _zz_shift_q_5 = shift_q_map_55;
      6'b111000 : _zz_shift_q_5 = shift_q_map_56;
      6'b111001 : _zz_shift_q_5 = shift_q_map_57;
      6'b111010 : _zz_shift_q_5 = shift_q_map_58;
      6'b111011 : _zz_shift_q_5 = shift_q_map_59;
      6'b111100 : _zz_shift_q_5 = shift_q_map_60;
      6'b111101 : _zz_shift_q_5 = shift_q_map_61;
      6'b111110 : _zz_shift_q_5 = shift_q_map_62;
      default : _zz_shift_q_5 = shift_q_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_6_1)
      6'b000000 : _zz_shift_i_6 = shift_i_map_0;
      6'b000001 : _zz_shift_i_6 = shift_i_map_1;
      6'b000010 : _zz_shift_i_6 = shift_i_map_2;
      6'b000011 : _zz_shift_i_6 = shift_i_map_3;
      6'b000100 : _zz_shift_i_6 = shift_i_map_4;
      6'b000101 : _zz_shift_i_6 = shift_i_map_5;
      6'b000110 : _zz_shift_i_6 = shift_i_map_6;
      6'b000111 : _zz_shift_i_6 = shift_i_map_7;
      6'b001000 : _zz_shift_i_6 = shift_i_map_8;
      6'b001001 : _zz_shift_i_6 = shift_i_map_9;
      6'b001010 : _zz_shift_i_6 = shift_i_map_10;
      6'b001011 : _zz_shift_i_6 = shift_i_map_11;
      6'b001100 : _zz_shift_i_6 = shift_i_map_12;
      6'b001101 : _zz_shift_i_6 = shift_i_map_13;
      6'b001110 : _zz_shift_i_6 = shift_i_map_14;
      6'b001111 : _zz_shift_i_6 = shift_i_map_15;
      6'b010000 : _zz_shift_i_6 = shift_i_map_16;
      6'b010001 : _zz_shift_i_6 = shift_i_map_17;
      6'b010010 : _zz_shift_i_6 = shift_i_map_18;
      6'b010011 : _zz_shift_i_6 = shift_i_map_19;
      6'b010100 : _zz_shift_i_6 = shift_i_map_20;
      6'b010101 : _zz_shift_i_6 = shift_i_map_21;
      6'b010110 : _zz_shift_i_6 = shift_i_map_22;
      6'b010111 : _zz_shift_i_6 = shift_i_map_23;
      6'b011000 : _zz_shift_i_6 = shift_i_map_24;
      6'b011001 : _zz_shift_i_6 = shift_i_map_25;
      6'b011010 : _zz_shift_i_6 = shift_i_map_26;
      6'b011011 : _zz_shift_i_6 = shift_i_map_27;
      6'b011100 : _zz_shift_i_6 = shift_i_map_28;
      6'b011101 : _zz_shift_i_6 = shift_i_map_29;
      6'b011110 : _zz_shift_i_6 = shift_i_map_30;
      6'b011111 : _zz_shift_i_6 = shift_i_map_31;
      6'b100000 : _zz_shift_i_6 = shift_i_map_32;
      6'b100001 : _zz_shift_i_6 = shift_i_map_33;
      6'b100010 : _zz_shift_i_6 = shift_i_map_34;
      6'b100011 : _zz_shift_i_6 = shift_i_map_35;
      6'b100100 : _zz_shift_i_6 = shift_i_map_36;
      6'b100101 : _zz_shift_i_6 = shift_i_map_37;
      6'b100110 : _zz_shift_i_6 = shift_i_map_38;
      6'b100111 : _zz_shift_i_6 = shift_i_map_39;
      6'b101000 : _zz_shift_i_6 = shift_i_map_40;
      6'b101001 : _zz_shift_i_6 = shift_i_map_41;
      6'b101010 : _zz_shift_i_6 = shift_i_map_42;
      6'b101011 : _zz_shift_i_6 = shift_i_map_43;
      6'b101100 : _zz_shift_i_6 = shift_i_map_44;
      6'b101101 : _zz_shift_i_6 = shift_i_map_45;
      6'b101110 : _zz_shift_i_6 = shift_i_map_46;
      6'b101111 : _zz_shift_i_6 = shift_i_map_47;
      6'b110000 : _zz_shift_i_6 = shift_i_map_48;
      6'b110001 : _zz_shift_i_6 = shift_i_map_49;
      6'b110010 : _zz_shift_i_6 = shift_i_map_50;
      6'b110011 : _zz_shift_i_6 = shift_i_map_51;
      6'b110100 : _zz_shift_i_6 = shift_i_map_52;
      6'b110101 : _zz_shift_i_6 = shift_i_map_53;
      6'b110110 : _zz_shift_i_6 = shift_i_map_54;
      6'b110111 : _zz_shift_i_6 = shift_i_map_55;
      6'b111000 : _zz_shift_i_6 = shift_i_map_56;
      6'b111001 : _zz_shift_i_6 = shift_i_map_57;
      6'b111010 : _zz_shift_i_6 = shift_i_map_58;
      6'b111011 : _zz_shift_i_6 = shift_i_map_59;
      6'b111100 : _zz_shift_i_6 = shift_i_map_60;
      6'b111101 : _zz_shift_i_6 = shift_i_map_61;
      6'b111110 : _zz_shift_i_6 = shift_i_map_62;
      default : _zz_shift_i_6 = shift_i_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_6_1)
      6'b000000 : _zz_shift_q_6 = shift_q_map_0;
      6'b000001 : _zz_shift_q_6 = shift_q_map_1;
      6'b000010 : _zz_shift_q_6 = shift_q_map_2;
      6'b000011 : _zz_shift_q_6 = shift_q_map_3;
      6'b000100 : _zz_shift_q_6 = shift_q_map_4;
      6'b000101 : _zz_shift_q_6 = shift_q_map_5;
      6'b000110 : _zz_shift_q_6 = shift_q_map_6;
      6'b000111 : _zz_shift_q_6 = shift_q_map_7;
      6'b001000 : _zz_shift_q_6 = shift_q_map_8;
      6'b001001 : _zz_shift_q_6 = shift_q_map_9;
      6'b001010 : _zz_shift_q_6 = shift_q_map_10;
      6'b001011 : _zz_shift_q_6 = shift_q_map_11;
      6'b001100 : _zz_shift_q_6 = shift_q_map_12;
      6'b001101 : _zz_shift_q_6 = shift_q_map_13;
      6'b001110 : _zz_shift_q_6 = shift_q_map_14;
      6'b001111 : _zz_shift_q_6 = shift_q_map_15;
      6'b010000 : _zz_shift_q_6 = shift_q_map_16;
      6'b010001 : _zz_shift_q_6 = shift_q_map_17;
      6'b010010 : _zz_shift_q_6 = shift_q_map_18;
      6'b010011 : _zz_shift_q_6 = shift_q_map_19;
      6'b010100 : _zz_shift_q_6 = shift_q_map_20;
      6'b010101 : _zz_shift_q_6 = shift_q_map_21;
      6'b010110 : _zz_shift_q_6 = shift_q_map_22;
      6'b010111 : _zz_shift_q_6 = shift_q_map_23;
      6'b011000 : _zz_shift_q_6 = shift_q_map_24;
      6'b011001 : _zz_shift_q_6 = shift_q_map_25;
      6'b011010 : _zz_shift_q_6 = shift_q_map_26;
      6'b011011 : _zz_shift_q_6 = shift_q_map_27;
      6'b011100 : _zz_shift_q_6 = shift_q_map_28;
      6'b011101 : _zz_shift_q_6 = shift_q_map_29;
      6'b011110 : _zz_shift_q_6 = shift_q_map_30;
      6'b011111 : _zz_shift_q_6 = shift_q_map_31;
      6'b100000 : _zz_shift_q_6 = shift_q_map_32;
      6'b100001 : _zz_shift_q_6 = shift_q_map_33;
      6'b100010 : _zz_shift_q_6 = shift_q_map_34;
      6'b100011 : _zz_shift_q_6 = shift_q_map_35;
      6'b100100 : _zz_shift_q_6 = shift_q_map_36;
      6'b100101 : _zz_shift_q_6 = shift_q_map_37;
      6'b100110 : _zz_shift_q_6 = shift_q_map_38;
      6'b100111 : _zz_shift_q_6 = shift_q_map_39;
      6'b101000 : _zz_shift_q_6 = shift_q_map_40;
      6'b101001 : _zz_shift_q_6 = shift_q_map_41;
      6'b101010 : _zz_shift_q_6 = shift_q_map_42;
      6'b101011 : _zz_shift_q_6 = shift_q_map_43;
      6'b101100 : _zz_shift_q_6 = shift_q_map_44;
      6'b101101 : _zz_shift_q_6 = shift_q_map_45;
      6'b101110 : _zz_shift_q_6 = shift_q_map_46;
      6'b101111 : _zz_shift_q_6 = shift_q_map_47;
      6'b110000 : _zz_shift_q_6 = shift_q_map_48;
      6'b110001 : _zz_shift_q_6 = shift_q_map_49;
      6'b110010 : _zz_shift_q_6 = shift_q_map_50;
      6'b110011 : _zz_shift_q_6 = shift_q_map_51;
      6'b110100 : _zz_shift_q_6 = shift_q_map_52;
      6'b110101 : _zz_shift_q_6 = shift_q_map_53;
      6'b110110 : _zz_shift_q_6 = shift_q_map_54;
      6'b110111 : _zz_shift_q_6 = shift_q_map_55;
      6'b111000 : _zz_shift_q_6 = shift_q_map_56;
      6'b111001 : _zz_shift_q_6 = shift_q_map_57;
      6'b111010 : _zz_shift_q_6 = shift_q_map_58;
      6'b111011 : _zz_shift_q_6 = shift_q_map_59;
      6'b111100 : _zz_shift_q_6 = shift_q_map_60;
      6'b111101 : _zz_shift_q_6 = shift_q_map_61;
      6'b111110 : _zz_shift_q_6 = shift_q_map_62;
      default : _zz_shift_q_6 = shift_q_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_7_1)
      6'b000000 : _zz_shift_i_7 = shift_i_map_0;
      6'b000001 : _zz_shift_i_7 = shift_i_map_1;
      6'b000010 : _zz_shift_i_7 = shift_i_map_2;
      6'b000011 : _zz_shift_i_7 = shift_i_map_3;
      6'b000100 : _zz_shift_i_7 = shift_i_map_4;
      6'b000101 : _zz_shift_i_7 = shift_i_map_5;
      6'b000110 : _zz_shift_i_7 = shift_i_map_6;
      6'b000111 : _zz_shift_i_7 = shift_i_map_7;
      6'b001000 : _zz_shift_i_7 = shift_i_map_8;
      6'b001001 : _zz_shift_i_7 = shift_i_map_9;
      6'b001010 : _zz_shift_i_7 = shift_i_map_10;
      6'b001011 : _zz_shift_i_7 = shift_i_map_11;
      6'b001100 : _zz_shift_i_7 = shift_i_map_12;
      6'b001101 : _zz_shift_i_7 = shift_i_map_13;
      6'b001110 : _zz_shift_i_7 = shift_i_map_14;
      6'b001111 : _zz_shift_i_7 = shift_i_map_15;
      6'b010000 : _zz_shift_i_7 = shift_i_map_16;
      6'b010001 : _zz_shift_i_7 = shift_i_map_17;
      6'b010010 : _zz_shift_i_7 = shift_i_map_18;
      6'b010011 : _zz_shift_i_7 = shift_i_map_19;
      6'b010100 : _zz_shift_i_7 = shift_i_map_20;
      6'b010101 : _zz_shift_i_7 = shift_i_map_21;
      6'b010110 : _zz_shift_i_7 = shift_i_map_22;
      6'b010111 : _zz_shift_i_7 = shift_i_map_23;
      6'b011000 : _zz_shift_i_7 = shift_i_map_24;
      6'b011001 : _zz_shift_i_7 = shift_i_map_25;
      6'b011010 : _zz_shift_i_7 = shift_i_map_26;
      6'b011011 : _zz_shift_i_7 = shift_i_map_27;
      6'b011100 : _zz_shift_i_7 = shift_i_map_28;
      6'b011101 : _zz_shift_i_7 = shift_i_map_29;
      6'b011110 : _zz_shift_i_7 = shift_i_map_30;
      6'b011111 : _zz_shift_i_7 = shift_i_map_31;
      6'b100000 : _zz_shift_i_7 = shift_i_map_32;
      6'b100001 : _zz_shift_i_7 = shift_i_map_33;
      6'b100010 : _zz_shift_i_7 = shift_i_map_34;
      6'b100011 : _zz_shift_i_7 = shift_i_map_35;
      6'b100100 : _zz_shift_i_7 = shift_i_map_36;
      6'b100101 : _zz_shift_i_7 = shift_i_map_37;
      6'b100110 : _zz_shift_i_7 = shift_i_map_38;
      6'b100111 : _zz_shift_i_7 = shift_i_map_39;
      6'b101000 : _zz_shift_i_7 = shift_i_map_40;
      6'b101001 : _zz_shift_i_7 = shift_i_map_41;
      6'b101010 : _zz_shift_i_7 = shift_i_map_42;
      6'b101011 : _zz_shift_i_7 = shift_i_map_43;
      6'b101100 : _zz_shift_i_7 = shift_i_map_44;
      6'b101101 : _zz_shift_i_7 = shift_i_map_45;
      6'b101110 : _zz_shift_i_7 = shift_i_map_46;
      6'b101111 : _zz_shift_i_7 = shift_i_map_47;
      6'b110000 : _zz_shift_i_7 = shift_i_map_48;
      6'b110001 : _zz_shift_i_7 = shift_i_map_49;
      6'b110010 : _zz_shift_i_7 = shift_i_map_50;
      6'b110011 : _zz_shift_i_7 = shift_i_map_51;
      6'b110100 : _zz_shift_i_7 = shift_i_map_52;
      6'b110101 : _zz_shift_i_7 = shift_i_map_53;
      6'b110110 : _zz_shift_i_7 = shift_i_map_54;
      6'b110111 : _zz_shift_i_7 = shift_i_map_55;
      6'b111000 : _zz_shift_i_7 = shift_i_map_56;
      6'b111001 : _zz_shift_i_7 = shift_i_map_57;
      6'b111010 : _zz_shift_i_7 = shift_i_map_58;
      6'b111011 : _zz_shift_i_7 = shift_i_map_59;
      6'b111100 : _zz_shift_i_7 = shift_i_map_60;
      6'b111101 : _zz_shift_i_7 = shift_i_map_61;
      6'b111110 : _zz_shift_i_7 = shift_i_map_62;
      default : _zz_shift_i_7 = shift_i_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_7_1)
      6'b000000 : _zz_shift_q_7 = shift_q_map_0;
      6'b000001 : _zz_shift_q_7 = shift_q_map_1;
      6'b000010 : _zz_shift_q_7 = shift_q_map_2;
      6'b000011 : _zz_shift_q_7 = shift_q_map_3;
      6'b000100 : _zz_shift_q_7 = shift_q_map_4;
      6'b000101 : _zz_shift_q_7 = shift_q_map_5;
      6'b000110 : _zz_shift_q_7 = shift_q_map_6;
      6'b000111 : _zz_shift_q_7 = shift_q_map_7;
      6'b001000 : _zz_shift_q_7 = shift_q_map_8;
      6'b001001 : _zz_shift_q_7 = shift_q_map_9;
      6'b001010 : _zz_shift_q_7 = shift_q_map_10;
      6'b001011 : _zz_shift_q_7 = shift_q_map_11;
      6'b001100 : _zz_shift_q_7 = shift_q_map_12;
      6'b001101 : _zz_shift_q_7 = shift_q_map_13;
      6'b001110 : _zz_shift_q_7 = shift_q_map_14;
      6'b001111 : _zz_shift_q_7 = shift_q_map_15;
      6'b010000 : _zz_shift_q_7 = shift_q_map_16;
      6'b010001 : _zz_shift_q_7 = shift_q_map_17;
      6'b010010 : _zz_shift_q_7 = shift_q_map_18;
      6'b010011 : _zz_shift_q_7 = shift_q_map_19;
      6'b010100 : _zz_shift_q_7 = shift_q_map_20;
      6'b010101 : _zz_shift_q_7 = shift_q_map_21;
      6'b010110 : _zz_shift_q_7 = shift_q_map_22;
      6'b010111 : _zz_shift_q_7 = shift_q_map_23;
      6'b011000 : _zz_shift_q_7 = shift_q_map_24;
      6'b011001 : _zz_shift_q_7 = shift_q_map_25;
      6'b011010 : _zz_shift_q_7 = shift_q_map_26;
      6'b011011 : _zz_shift_q_7 = shift_q_map_27;
      6'b011100 : _zz_shift_q_7 = shift_q_map_28;
      6'b011101 : _zz_shift_q_7 = shift_q_map_29;
      6'b011110 : _zz_shift_q_7 = shift_q_map_30;
      6'b011111 : _zz_shift_q_7 = shift_q_map_31;
      6'b100000 : _zz_shift_q_7 = shift_q_map_32;
      6'b100001 : _zz_shift_q_7 = shift_q_map_33;
      6'b100010 : _zz_shift_q_7 = shift_q_map_34;
      6'b100011 : _zz_shift_q_7 = shift_q_map_35;
      6'b100100 : _zz_shift_q_7 = shift_q_map_36;
      6'b100101 : _zz_shift_q_7 = shift_q_map_37;
      6'b100110 : _zz_shift_q_7 = shift_q_map_38;
      6'b100111 : _zz_shift_q_7 = shift_q_map_39;
      6'b101000 : _zz_shift_q_7 = shift_q_map_40;
      6'b101001 : _zz_shift_q_7 = shift_q_map_41;
      6'b101010 : _zz_shift_q_7 = shift_q_map_42;
      6'b101011 : _zz_shift_q_7 = shift_q_map_43;
      6'b101100 : _zz_shift_q_7 = shift_q_map_44;
      6'b101101 : _zz_shift_q_7 = shift_q_map_45;
      6'b101110 : _zz_shift_q_7 = shift_q_map_46;
      6'b101111 : _zz_shift_q_7 = shift_q_map_47;
      6'b110000 : _zz_shift_q_7 = shift_q_map_48;
      6'b110001 : _zz_shift_q_7 = shift_q_map_49;
      6'b110010 : _zz_shift_q_7 = shift_q_map_50;
      6'b110011 : _zz_shift_q_7 = shift_q_map_51;
      6'b110100 : _zz_shift_q_7 = shift_q_map_52;
      6'b110101 : _zz_shift_q_7 = shift_q_map_53;
      6'b110110 : _zz_shift_q_7 = shift_q_map_54;
      6'b110111 : _zz_shift_q_7 = shift_q_map_55;
      6'b111000 : _zz_shift_q_7 = shift_q_map_56;
      6'b111001 : _zz_shift_q_7 = shift_q_map_57;
      6'b111010 : _zz_shift_q_7 = shift_q_map_58;
      6'b111011 : _zz_shift_q_7 = shift_q_map_59;
      6'b111100 : _zz_shift_q_7 = shift_q_map_60;
      6'b111101 : _zz_shift_q_7 = shift_q_map_61;
      6'b111110 : _zz_shift_q_7 = shift_q_map_62;
      default : _zz_shift_q_7 = shift_q_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_0_3)
      6'b000000 : _zz_shift_i_0_2 = shift_i_map_0;
      6'b000001 : _zz_shift_i_0_2 = shift_i_map_1;
      6'b000010 : _zz_shift_i_0_2 = shift_i_map_2;
      6'b000011 : _zz_shift_i_0_2 = shift_i_map_3;
      6'b000100 : _zz_shift_i_0_2 = shift_i_map_4;
      6'b000101 : _zz_shift_i_0_2 = shift_i_map_5;
      6'b000110 : _zz_shift_i_0_2 = shift_i_map_6;
      6'b000111 : _zz_shift_i_0_2 = shift_i_map_7;
      6'b001000 : _zz_shift_i_0_2 = shift_i_map_8;
      6'b001001 : _zz_shift_i_0_2 = shift_i_map_9;
      6'b001010 : _zz_shift_i_0_2 = shift_i_map_10;
      6'b001011 : _zz_shift_i_0_2 = shift_i_map_11;
      6'b001100 : _zz_shift_i_0_2 = shift_i_map_12;
      6'b001101 : _zz_shift_i_0_2 = shift_i_map_13;
      6'b001110 : _zz_shift_i_0_2 = shift_i_map_14;
      6'b001111 : _zz_shift_i_0_2 = shift_i_map_15;
      6'b010000 : _zz_shift_i_0_2 = shift_i_map_16;
      6'b010001 : _zz_shift_i_0_2 = shift_i_map_17;
      6'b010010 : _zz_shift_i_0_2 = shift_i_map_18;
      6'b010011 : _zz_shift_i_0_2 = shift_i_map_19;
      6'b010100 : _zz_shift_i_0_2 = shift_i_map_20;
      6'b010101 : _zz_shift_i_0_2 = shift_i_map_21;
      6'b010110 : _zz_shift_i_0_2 = shift_i_map_22;
      6'b010111 : _zz_shift_i_0_2 = shift_i_map_23;
      6'b011000 : _zz_shift_i_0_2 = shift_i_map_24;
      6'b011001 : _zz_shift_i_0_2 = shift_i_map_25;
      6'b011010 : _zz_shift_i_0_2 = shift_i_map_26;
      6'b011011 : _zz_shift_i_0_2 = shift_i_map_27;
      6'b011100 : _zz_shift_i_0_2 = shift_i_map_28;
      6'b011101 : _zz_shift_i_0_2 = shift_i_map_29;
      6'b011110 : _zz_shift_i_0_2 = shift_i_map_30;
      6'b011111 : _zz_shift_i_0_2 = shift_i_map_31;
      6'b100000 : _zz_shift_i_0_2 = shift_i_map_32;
      6'b100001 : _zz_shift_i_0_2 = shift_i_map_33;
      6'b100010 : _zz_shift_i_0_2 = shift_i_map_34;
      6'b100011 : _zz_shift_i_0_2 = shift_i_map_35;
      6'b100100 : _zz_shift_i_0_2 = shift_i_map_36;
      6'b100101 : _zz_shift_i_0_2 = shift_i_map_37;
      6'b100110 : _zz_shift_i_0_2 = shift_i_map_38;
      6'b100111 : _zz_shift_i_0_2 = shift_i_map_39;
      6'b101000 : _zz_shift_i_0_2 = shift_i_map_40;
      6'b101001 : _zz_shift_i_0_2 = shift_i_map_41;
      6'b101010 : _zz_shift_i_0_2 = shift_i_map_42;
      6'b101011 : _zz_shift_i_0_2 = shift_i_map_43;
      6'b101100 : _zz_shift_i_0_2 = shift_i_map_44;
      6'b101101 : _zz_shift_i_0_2 = shift_i_map_45;
      6'b101110 : _zz_shift_i_0_2 = shift_i_map_46;
      6'b101111 : _zz_shift_i_0_2 = shift_i_map_47;
      6'b110000 : _zz_shift_i_0_2 = shift_i_map_48;
      6'b110001 : _zz_shift_i_0_2 = shift_i_map_49;
      6'b110010 : _zz_shift_i_0_2 = shift_i_map_50;
      6'b110011 : _zz_shift_i_0_2 = shift_i_map_51;
      6'b110100 : _zz_shift_i_0_2 = shift_i_map_52;
      6'b110101 : _zz_shift_i_0_2 = shift_i_map_53;
      6'b110110 : _zz_shift_i_0_2 = shift_i_map_54;
      6'b110111 : _zz_shift_i_0_2 = shift_i_map_55;
      6'b111000 : _zz_shift_i_0_2 = shift_i_map_56;
      6'b111001 : _zz_shift_i_0_2 = shift_i_map_57;
      6'b111010 : _zz_shift_i_0_2 = shift_i_map_58;
      6'b111011 : _zz_shift_i_0_2 = shift_i_map_59;
      6'b111100 : _zz_shift_i_0_2 = shift_i_map_60;
      6'b111101 : _zz_shift_i_0_2 = shift_i_map_61;
      6'b111110 : _zz_shift_i_0_2 = shift_i_map_62;
      default : _zz_shift_i_0_2 = shift_i_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_0_3)
      6'b000000 : _zz_shift_q_0_2 = shift_q_map_0;
      6'b000001 : _zz_shift_q_0_2 = shift_q_map_1;
      6'b000010 : _zz_shift_q_0_2 = shift_q_map_2;
      6'b000011 : _zz_shift_q_0_2 = shift_q_map_3;
      6'b000100 : _zz_shift_q_0_2 = shift_q_map_4;
      6'b000101 : _zz_shift_q_0_2 = shift_q_map_5;
      6'b000110 : _zz_shift_q_0_2 = shift_q_map_6;
      6'b000111 : _zz_shift_q_0_2 = shift_q_map_7;
      6'b001000 : _zz_shift_q_0_2 = shift_q_map_8;
      6'b001001 : _zz_shift_q_0_2 = shift_q_map_9;
      6'b001010 : _zz_shift_q_0_2 = shift_q_map_10;
      6'b001011 : _zz_shift_q_0_2 = shift_q_map_11;
      6'b001100 : _zz_shift_q_0_2 = shift_q_map_12;
      6'b001101 : _zz_shift_q_0_2 = shift_q_map_13;
      6'b001110 : _zz_shift_q_0_2 = shift_q_map_14;
      6'b001111 : _zz_shift_q_0_2 = shift_q_map_15;
      6'b010000 : _zz_shift_q_0_2 = shift_q_map_16;
      6'b010001 : _zz_shift_q_0_2 = shift_q_map_17;
      6'b010010 : _zz_shift_q_0_2 = shift_q_map_18;
      6'b010011 : _zz_shift_q_0_2 = shift_q_map_19;
      6'b010100 : _zz_shift_q_0_2 = shift_q_map_20;
      6'b010101 : _zz_shift_q_0_2 = shift_q_map_21;
      6'b010110 : _zz_shift_q_0_2 = shift_q_map_22;
      6'b010111 : _zz_shift_q_0_2 = shift_q_map_23;
      6'b011000 : _zz_shift_q_0_2 = shift_q_map_24;
      6'b011001 : _zz_shift_q_0_2 = shift_q_map_25;
      6'b011010 : _zz_shift_q_0_2 = shift_q_map_26;
      6'b011011 : _zz_shift_q_0_2 = shift_q_map_27;
      6'b011100 : _zz_shift_q_0_2 = shift_q_map_28;
      6'b011101 : _zz_shift_q_0_2 = shift_q_map_29;
      6'b011110 : _zz_shift_q_0_2 = shift_q_map_30;
      6'b011111 : _zz_shift_q_0_2 = shift_q_map_31;
      6'b100000 : _zz_shift_q_0_2 = shift_q_map_32;
      6'b100001 : _zz_shift_q_0_2 = shift_q_map_33;
      6'b100010 : _zz_shift_q_0_2 = shift_q_map_34;
      6'b100011 : _zz_shift_q_0_2 = shift_q_map_35;
      6'b100100 : _zz_shift_q_0_2 = shift_q_map_36;
      6'b100101 : _zz_shift_q_0_2 = shift_q_map_37;
      6'b100110 : _zz_shift_q_0_2 = shift_q_map_38;
      6'b100111 : _zz_shift_q_0_2 = shift_q_map_39;
      6'b101000 : _zz_shift_q_0_2 = shift_q_map_40;
      6'b101001 : _zz_shift_q_0_2 = shift_q_map_41;
      6'b101010 : _zz_shift_q_0_2 = shift_q_map_42;
      6'b101011 : _zz_shift_q_0_2 = shift_q_map_43;
      6'b101100 : _zz_shift_q_0_2 = shift_q_map_44;
      6'b101101 : _zz_shift_q_0_2 = shift_q_map_45;
      6'b101110 : _zz_shift_q_0_2 = shift_q_map_46;
      6'b101111 : _zz_shift_q_0_2 = shift_q_map_47;
      6'b110000 : _zz_shift_q_0_2 = shift_q_map_48;
      6'b110001 : _zz_shift_q_0_2 = shift_q_map_49;
      6'b110010 : _zz_shift_q_0_2 = shift_q_map_50;
      6'b110011 : _zz_shift_q_0_2 = shift_q_map_51;
      6'b110100 : _zz_shift_q_0_2 = shift_q_map_52;
      6'b110101 : _zz_shift_q_0_2 = shift_q_map_53;
      6'b110110 : _zz_shift_q_0_2 = shift_q_map_54;
      6'b110111 : _zz_shift_q_0_2 = shift_q_map_55;
      6'b111000 : _zz_shift_q_0_2 = shift_q_map_56;
      6'b111001 : _zz_shift_q_0_2 = shift_q_map_57;
      6'b111010 : _zz_shift_q_0_2 = shift_q_map_58;
      6'b111011 : _zz_shift_q_0_2 = shift_q_map_59;
      6'b111100 : _zz_shift_q_0_2 = shift_q_map_60;
      6'b111101 : _zz_shift_q_0_2 = shift_q_map_61;
      6'b111110 : _zz_shift_q_0_2 = shift_q_map_62;
      default : _zz_shift_q_0_2 = shift_q_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_1_3)
      6'b000000 : _zz_shift_i_1_2 = shift_i_map_0;
      6'b000001 : _zz_shift_i_1_2 = shift_i_map_1;
      6'b000010 : _zz_shift_i_1_2 = shift_i_map_2;
      6'b000011 : _zz_shift_i_1_2 = shift_i_map_3;
      6'b000100 : _zz_shift_i_1_2 = shift_i_map_4;
      6'b000101 : _zz_shift_i_1_2 = shift_i_map_5;
      6'b000110 : _zz_shift_i_1_2 = shift_i_map_6;
      6'b000111 : _zz_shift_i_1_2 = shift_i_map_7;
      6'b001000 : _zz_shift_i_1_2 = shift_i_map_8;
      6'b001001 : _zz_shift_i_1_2 = shift_i_map_9;
      6'b001010 : _zz_shift_i_1_2 = shift_i_map_10;
      6'b001011 : _zz_shift_i_1_2 = shift_i_map_11;
      6'b001100 : _zz_shift_i_1_2 = shift_i_map_12;
      6'b001101 : _zz_shift_i_1_2 = shift_i_map_13;
      6'b001110 : _zz_shift_i_1_2 = shift_i_map_14;
      6'b001111 : _zz_shift_i_1_2 = shift_i_map_15;
      6'b010000 : _zz_shift_i_1_2 = shift_i_map_16;
      6'b010001 : _zz_shift_i_1_2 = shift_i_map_17;
      6'b010010 : _zz_shift_i_1_2 = shift_i_map_18;
      6'b010011 : _zz_shift_i_1_2 = shift_i_map_19;
      6'b010100 : _zz_shift_i_1_2 = shift_i_map_20;
      6'b010101 : _zz_shift_i_1_2 = shift_i_map_21;
      6'b010110 : _zz_shift_i_1_2 = shift_i_map_22;
      6'b010111 : _zz_shift_i_1_2 = shift_i_map_23;
      6'b011000 : _zz_shift_i_1_2 = shift_i_map_24;
      6'b011001 : _zz_shift_i_1_2 = shift_i_map_25;
      6'b011010 : _zz_shift_i_1_2 = shift_i_map_26;
      6'b011011 : _zz_shift_i_1_2 = shift_i_map_27;
      6'b011100 : _zz_shift_i_1_2 = shift_i_map_28;
      6'b011101 : _zz_shift_i_1_2 = shift_i_map_29;
      6'b011110 : _zz_shift_i_1_2 = shift_i_map_30;
      6'b011111 : _zz_shift_i_1_2 = shift_i_map_31;
      6'b100000 : _zz_shift_i_1_2 = shift_i_map_32;
      6'b100001 : _zz_shift_i_1_2 = shift_i_map_33;
      6'b100010 : _zz_shift_i_1_2 = shift_i_map_34;
      6'b100011 : _zz_shift_i_1_2 = shift_i_map_35;
      6'b100100 : _zz_shift_i_1_2 = shift_i_map_36;
      6'b100101 : _zz_shift_i_1_2 = shift_i_map_37;
      6'b100110 : _zz_shift_i_1_2 = shift_i_map_38;
      6'b100111 : _zz_shift_i_1_2 = shift_i_map_39;
      6'b101000 : _zz_shift_i_1_2 = shift_i_map_40;
      6'b101001 : _zz_shift_i_1_2 = shift_i_map_41;
      6'b101010 : _zz_shift_i_1_2 = shift_i_map_42;
      6'b101011 : _zz_shift_i_1_2 = shift_i_map_43;
      6'b101100 : _zz_shift_i_1_2 = shift_i_map_44;
      6'b101101 : _zz_shift_i_1_2 = shift_i_map_45;
      6'b101110 : _zz_shift_i_1_2 = shift_i_map_46;
      6'b101111 : _zz_shift_i_1_2 = shift_i_map_47;
      6'b110000 : _zz_shift_i_1_2 = shift_i_map_48;
      6'b110001 : _zz_shift_i_1_2 = shift_i_map_49;
      6'b110010 : _zz_shift_i_1_2 = shift_i_map_50;
      6'b110011 : _zz_shift_i_1_2 = shift_i_map_51;
      6'b110100 : _zz_shift_i_1_2 = shift_i_map_52;
      6'b110101 : _zz_shift_i_1_2 = shift_i_map_53;
      6'b110110 : _zz_shift_i_1_2 = shift_i_map_54;
      6'b110111 : _zz_shift_i_1_2 = shift_i_map_55;
      6'b111000 : _zz_shift_i_1_2 = shift_i_map_56;
      6'b111001 : _zz_shift_i_1_2 = shift_i_map_57;
      6'b111010 : _zz_shift_i_1_2 = shift_i_map_58;
      6'b111011 : _zz_shift_i_1_2 = shift_i_map_59;
      6'b111100 : _zz_shift_i_1_2 = shift_i_map_60;
      6'b111101 : _zz_shift_i_1_2 = shift_i_map_61;
      6'b111110 : _zz_shift_i_1_2 = shift_i_map_62;
      default : _zz_shift_i_1_2 = shift_i_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_1_3)
      6'b000000 : _zz_shift_q_1_2 = shift_q_map_0;
      6'b000001 : _zz_shift_q_1_2 = shift_q_map_1;
      6'b000010 : _zz_shift_q_1_2 = shift_q_map_2;
      6'b000011 : _zz_shift_q_1_2 = shift_q_map_3;
      6'b000100 : _zz_shift_q_1_2 = shift_q_map_4;
      6'b000101 : _zz_shift_q_1_2 = shift_q_map_5;
      6'b000110 : _zz_shift_q_1_2 = shift_q_map_6;
      6'b000111 : _zz_shift_q_1_2 = shift_q_map_7;
      6'b001000 : _zz_shift_q_1_2 = shift_q_map_8;
      6'b001001 : _zz_shift_q_1_2 = shift_q_map_9;
      6'b001010 : _zz_shift_q_1_2 = shift_q_map_10;
      6'b001011 : _zz_shift_q_1_2 = shift_q_map_11;
      6'b001100 : _zz_shift_q_1_2 = shift_q_map_12;
      6'b001101 : _zz_shift_q_1_2 = shift_q_map_13;
      6'b001110 : _zz_shift_q_1_2 = shift_q_map_14;
      6'b001111 : _zz_shift_q_1_2 = shift_q_map_15;
      6'b010000 : _zz_shift_q_1_2 = shift_q_map_16;
      6'b010001 : _zz_shift_q_1_2 = shift_q_map_17;
      6'b010010 : _zz_shift_q_1_2 = shift_q_map_18;
      6'b010011 : _zz_shift_q_1_2 = shift_q_map_19;
      6'b010100 : _zz_shift_q_1_2 = shift_q_map_20;
      6'b010101 : _zz_shift_q_1_2 = shift_q_map_21;
      6'b010110 : _zz_shift_q_1_2 = shift_q_map_22;
      6'b010111 : _zz_shift_q_1_2 = shift_q_map_23;
      6'b011000 : _zz_shift_q_1_2 = shift_q_map_24;
      6'b011001 : _zz_shift_q_1_2 = shift_q_map_25;
      6'b011010 : _zz_shift_q_1_2 = shift_q_map_26;
      6'b011011 : _zz_shift_q_1_2 = shift_q_map_27;
      6'b011100 : _zz_shift_q_1_2 = shift_q_map_28;
      6'b011101 : _zz_shift_q_1_2 = shift_q_map_29;
      6'b011110 : _zz_shift_q_1_2 = shift_q_map_30;
      6'b011111 : _zz_shift_q_1_2 = shift_q_map_31;
      6'b100000 : _zz_shift_q_1_2 = shift_q_map_32;
      6'b100001 : _zz_shift_q_1_2 = shift_q_map_33;
      6'b100010 : _zz_shift_q_1_2 = shift_q_map_34;
      6'b100011 : _zz_shift_q_1_2 = shift_q_map_35;
      6'b100100 : _zz_shift_q_1_2 = shift_q_map_36;
      6'b100101 : _zz_shift_q_1_2 = shift_q_map_37;
      6'b100110 : _zz_shift_q_1_2 = shift_q_map_38;
      6'b100111 : _zz_shift_q_1_2 = shift_q_map_39;
      6'b101000 : _zz_shift_q_1_2 = shift_q_map_40;
      6'b101001 : _zz_shift_q_1_2 = shift_q_map_41;
      6'b101010 : _zz_shift_q_1_2 = shift_q_map_42;
      6'b101011 : _zz_shift_q_1_2 = shift_q_map_43;
      6'b101100 : _zz_shift_q_1_2 = shift_q_map_44;
      6'b101101 : _zz_shift_q_1_2 = shift_q_map_45;
      6'b101110 : _zz_shift_q_1_2 = shift_q_map_46;
      6'b101111 : _zz_shift_q_1_2 = shift_q_map_47;
      6'b110000 : _zz_shift_q_1_2 = shift_q_map_48;
      6'b110001 : _zz_shift_q_1_2 = shift_q_map_49;
      6'b110010 : _zz_shift_q_1_2 = shift_q_map_50;
      6'b110011 : _zz_shift_q_1_2 = shift_q_map_51;
      6'b110100 : _zz_shift_q_1_2 = shift_q_map_52;
      6'b110101 : _zz_shift_q_1_2 = shift_q_map_53;
      6'b110110 : _zz_shift_q_1_2 = shift_q_map_54;
      6'b110111 : _zz_shift_q_1_2 = shift_q_map_55;
      6'b111000 : _zz_shift_q_1_2 = shift_q_map_56;
      6'b111001 : _zz_shift_q_1_2 = shift_q_map_57;
      6'b111010 : _zz_shift_q_1_2 = shift_q_map_58;
      6'b111011 : _zz_shift_q_1_2 = shift_q_map_59;
      6'b111100 : _zz_shift_q_1_2 = shift_q_map_60;
      6'b111101 : _zz_shift_q_1_2 = shift_q_map_61;
      6'b111110 : _zz_shift_q_1_2 = shift_q_map_62;
      default : _zz_shift_q_1_2 = shift_q_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_2_3)
      6'b000000 : _zz_shift_i_2_2 = shift_i_map_0;
      6'b000001 : _zz_shift_i_2_2 = shift_i_map_1;
      6'b000010 : _zz_shift_i_2_2 = shift_i_map_2;
      6'b000011 : _zz_shift_i_2_2 = shift_i_map_3;
      6'b000100 : _zz_shift_i_2_2 = shift_i_map_4;
      6'b000101 : _zz_shift_i_2_2 = shift_i_map_5;
      6'b000110 : _zz_shift_i_2_2 = shift_i_map_6;
      6'b000111 : _zz_shift_i_2_2 = shift_i_map_7;
      6'b001000 : _zz_shift_i_2_2 = shift_i_map_8;
      6'b001001 : _zz_shift_i_2_2 = shift_i_map_9;
      6'b001010 : _zz_shift_i_2_2 = shift_i_map_10;
      6'b001011 : _zz_shift_i_2_2 = shift_i_map_11;
      6'b001100 : _zz_shift_i_2_2 = shift_i_map_12;
      6'b001101 : _zz_shift_i_2_2 = shift_i_map_13;
      6'b001110 : _zz_shift_i_2_2 = shift_i_map_14;
      6'b001111 : _zz_shift_i_2_2 = shift_i_map_15;
      6'b010000 : _zz_shift_i_2_2 = shift_i_map_16;
      6'b010001 : _zz_shift_i_2_2 = shift_i_map_17;
      6'b010010 : _zz_shift_i_2_2 = shift_i_map_18;
      6'b010011 : _zz_shift_i_2_2 = shift_i_map_19;
      6'b010100 : _zz_shift_i_2_2 = shift_i_map_20;
      6'b010101 : _zz_shift_i_2_2 = shift_i_map_21;
      6'b010110 : _zz_shift_i_2_2 = shift_i_map_22;
      6'b010111 : _zz_shift_i_2_2 = shift_i_map_23;
      6'b011000 : _zz_shift_i_2_2 = shift_i_map_24;
      6'b011001 : _zz_shift_i_2_2 = shift_i_map_25;
      6'b011010 : _zz_shift_i_2_2 = shift_i_map_26;
      6'b011011 : _zz_shift_i_2_2 = shift_i_map_27;
      6'b011100 : _zz_shift_i_2_2 = shift_i_map_28;
      6'b011101 : _zz_shift_i_2_2 = shift_i_map_29;
      6'b011110 : _zz_shift_i_2_2 = shift_i_map_30;
      6'b011111 : _zz_shift_i_2_2 = shift_i_map_31;
      6'b100000 : _zz_shift_i_2_2 = shift_i_map_32;
      6'b100001 : _zz_shift_i_2_2 = shift_i_map_33;
      6'b100010 : _zz_shift_i_2_2 = shift_i_map_34;
      6'b100011 : _zz_shift_i_2_2 = shift_i_map_35;
      6'b100100 : _zz_shift_i_2_2 = shift_i_map_36;
      6'b100101 : _zz_shift_i_2_2 = shift_i_map_37;
      6'b100110 : _zz_shift_i_2_2 = shift_i_map_38;
      6'b100111 : _zz_shift_i_2_2 = shift_i_map_39;
      6'b101000 : _zz_shift_i_2_2 = shift_i_map_40;
      6'b101001 : _zz_shift_i_2_2 = shift_i_map_41;
      6'b101010 : _zz_shift_i_2_2 = shift_i_map_42;
      6'b101011 : _zz_shift_i_2_2 = shift_i_map_43;
      6'b101100 : _zz_shift_i_2_2 = shift_i_map_44;
      6'b101101 : _zz_shift_i_2_2 = shift_i_map_45;
      6'b101110 : _zz_shift_i_2_2 = shift_i_map_46;
      6'b101111 : _zz_shift_i_2_2 = shift_i_map_47;
      6'b110000 : _zz_shift_i_2_2 = shift_i_map_48;
      6'b110001 : _zz_shift_i_2_2 = shift_i_map_49;
      6'b110010 : _zz_shift_i_2_2 = shift_i_map_50;
      6'b110011 : _zz_shift_i_2_2 = shift_i_map_51;
      6'b110100 : _zz_shift_i_2_2 = shift_i_map_52;
      6'b110101 : _zz_shift_i_2_2 = shift_i_map_53;
      6'b110110 : _zz_shift_i_2_2 = shift_i_map_54;
      6'b110111 : _zz_shift_i_2_2 = shift_i_map_55;
      6'b111000 : _zz_shift_i_2_2 = shift_i_map_56;
      6'b111001 : _zz_shift_i_2_2 = shift_i_map_57;
      6'b111010 : _zz_shift_i_2_2 = shift_i_map_58;
      6'b111011 : _zz_shift_i_2_2 = shift_i_map_59;
      6'b111100 : _zz_shift_i_2_2 = shift_i_map_60;
      6'b111101 : _zz_shift_i_2_2 = shift_i_map_61;
      6'b111110 : _zz_shift_i_2_2 = shift_i_map_62;
      default : _zz_shift_i_2_2 = shift_i_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_2_3)
      6'b000000 : _zz_shift_q_2_2 = shift_q_map_0;
      6'b000001 : _zz_shift_q_2_2 = shift_q_map_1;
      6'b000010 : _zz_shift_q_2_2 = shift_q_map_2;
      6'b000011 : _zz_shift_q_2_2 = shift_q_map_3;
      6'b000100 : _zz_shift_q_2_2 = shift_q_map_4;
      6'b000101 : _zz_shift_q_2_2 = shift_q_map_5;
      6'b000110 : _zz_shift_q_2_2 = shift_q_map_6;
      6'b000111 : _zz_shift_q_2_2 = shift_q_map_7;
      6'b001000 : _zz_shift_q_2_2 = shift_q_map_8;
      6'b001001 : _zz_shift_q_2_2 = shift_q_map_9;
      6'b001010 : _zz_shift_q_2_2 = shift_q_map_10;
      6'b001011 : _zz_shift_q_2_2 = shift_q_map_11;
      6'b001100 : _zz_shift_q_2_2 = shift_q_map_12;
      6'b001101 : _zz_shift_q_2_2 = shift_q_map_13;
      6'b001110 : _zz_shift_q_2_2 = shift_q_map_14;
      6'b001111 : _zz_shift_q_2_2 = shift_q_map_15;
      6'b010000 : _zz_shift_q_2_2 = shift_q_map_16;
      6'b010001 : _zz_shift_q_2_2 = shift_q_map_17;
      6'b010010 : _zz_shift_q_2_2 = shift_q_map_18;
      6'b010011 : _zz_shift_q_2_2 = shift_q_map_19;
      6'b010100 : _zz_shift_q_2_2 = shift_q_map_20;
      6'b010101 : _zz_shift_q_2_2 = shift_q_map_21;
      6'b010110 : _zz_shift_q_2_2 = shift_q_map_22;
      6'b010111 : _zz_shift_q_2_2 = shift_q_map_23;
      6'b011000 : _zz_shift_q_2_2 = shift_q_map_24;
      6'b011001 : _zz_shift_q_2_2 = shift_q_map_25;
      6'b011010 : _zz_shift_q_2_2 = shift_q_map_26;
      6'b011011 : _zz_shift_q_2_2 = shift_q_map_27;
      6'b011100 : _zz_shift_q_2_2 = shift_q_map_28;
      6'b011101 : _zz_shift_q_2_2 = shift_q_map_29;
      6'b011110 : _zz_shift_q_2_2 = shift_q_map_30;
      6'b011111 : _zz_shift_q_2_2 = shift_q_map_31;
      6'b100000 : _zz_shift_q_2_2 = shift_q_map_32;
      6'b100001 : _zz_shift_q_2_2 = shift_q_map_33;
      6'b100010 : _zz_shift_q_2_2 = shift_q_map_34;
      6'b100011 : _zz_shift_q_2_2 = shift_q_map_35;
      6'b100100 : _zz_shift_q_2_2 = shift_q_map_36;
      6'b100101 : _zz_shift_q_2_2 = shift_q_map_37;
      6'b100110 : _zz_shift_q_2_2 = shift_q_map_38;
      6'b100111 : _zz_shift_q_2_2 = shift_q_map_39;
      6'b101000 : _zz_shift_q_2_2 = shift_q_map_40;
      6'b101001 : _zz_shift_q_2_2 = shift_q_map_41;
      6'b101010 : _zz_shift_q_2_2 = shift_q_map_42;
      6'b101011 : _zz_shift_q_2_2 = shift_q_map_43;
      6'b101100 : _zz_shift_q_2_2 = shift_q_map_44;
      6'b101101 : _zz_shift_q_2_2 = shift_q_map_45;
      6'b101110 : _zz_shift_q_2_2 = shift_q_map_46;
      6'b101111 : _zz_shift_q_2_2 = shift_q_map_47;
      6'b110000 : _zz_shift_q_2_2 = shift_q_map_48;
      6'b110001 : _zz_shift_q_2_2 = shift_q_map_49;
      6'b110010 : _zz_shift_q_2_2 = shift_q_map_50;
      6'b110011 : _zz_shift_q_2_2 = shift_q_map_51;
      6'b110100 : _zz_shift_q_2_2 = shift_q_map_52;
      6'b110101 : _zz_shift_q_2_2 = shift_q_map_53;
      6'b110110 : _zz_shift_q_2_2 = shift_q_map_54;
      6'b110111 : _zz_shift_q_2_2 = shift_q_map_55;
      6'b111000 : _zz_shift_q_2_2 = shift_q_map_56;
      6'b111001 : _zz_shift_q_2_2 = shift_q_map_57;
      6'b111010 : _zz_shift_q_2_2 = shift_q_map_58;
      6'b111011 : _zz_shift_q_2_2 = shift_q_map_59;
      6'b111100 : _zz_shift_q_2_2 = shift_q_map_60;
      6'b111101 : _zz_shift_q_2_2 = shift_q_map_61;
      6'b111110 : _zz_shift_q_2_2 = shift_q_map_62;
      default : _zz_shift_q_2_2 = shift_q_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_3_3)
      6'b000000 : _zz_shift_i_3_2 = shift_i_map_0;
      6'b000001 : _zz_shift_i_3_2 = shift_i_map_1;
      6'b000010 : _zz_shift_i_3_2 = shift_i_map_2;
      6'b000011 : _zz_shift_i_3_2 = shift_i_map_3;
      6'b000100 : _zz_shift_i_3_2 = shift_i_map_4;
      6'b000101 : _zz_shift_i_3_2 = shift_i_map_5;
      6'b000110 : _zz_shift_i_3_2 = shift_i_map_6;
      6'b000111 : _zz_shift_i_3_2 = shift_i_map_7;
      6'b001000 : _zz_shift_i_3_2 = shift_i_map_8;
      6'b001001 : _zz_shift_i_3_2 = shift_i_map_9;
      6'b001010 : _zz_shift_i_3_2 = shift_i_map_10;
      6'b001011 : _zz_shift_i_3_2 = shift_i_map_11;
      6'b001100 : _zz_shift_i_3_2 = shift_i_map_12;
      6'b001101 : _zz_shift_i_3_2 = shift_i_map_13;
      6'b001110 : _zz_shift_i_3_2 = shift_i_map_14;
      6'b001111 : _zz_shift_i_3_2 = shift_i_map_15;
      6'b010000 : _zz_shift_i_3_2 = shift_i_map_16;
      6'b010001 : _zz_shift_i_3_2 = shift_i_map_17;
      6'b010010 : _zz_shift_i_3_2 = shift_i_map_18;
      6'b010011 : _zz_shift_i_3_2 = shift_i_map_19;
      6'b010100 : _zz_shift_i_3_2 = shift_i_map_20;
      6'b010101 : _zz_shift_i_3_2 = shift_i_map_21;
      6'b010110 : _zz_shift_i_3_2 = shift_i_map_22;
      6'b010111 : _zz_shift_i_3_2 = shift_i_map_23;
      6'b011000 : _zz_shift_i_3_2 = shift_i_map_24;
      6'b011001 : _zz_shift_i_3_2 = shift_i_map_25;
      6'b011010 : _zz_shift_i_3_2 = shift_i_map_26;
      6'b011011 : _zz_shift_i_3_2 = shift_i_map_27;
      6'b011100 : _zz_shift_i_3_2 = shift_i_map_28;
      6'b011101 : _zz_shift_i_3_2 = shift_i_map_29;
      6'b011110 : _zz_shift_i_3_2 = shift_i_map_30;
      6'b011111 : _zz_shift_i_3_2 = shift_i_map_31;
      6'b100000 : _zz_shift_i_3_2 = shift_i_map_32;
      6'b100001 : _zz_shift_i_3_2 = shift_i_map_33;
      6'b100010 : _zz_shift_i_3_2 = shift_i_map_34;
      6'b100011 : _zz_shift_i_3_2 = shift_i_map_35;
      6'b100100 : _zz_shift_i_3_2 = shift_i_map_36;
      6'b100101 : _zz_shift_i_3_2 = shift_i_map_37;
      6'b100110 : _zz_shift_i_3_2 = shift_i_map_38;
      6'b100111 : _zz_shift_i_3_2 = shift_i_map_39;
      6'b101000 : _zz_shift_i_3_2 = shift_i_map_40;
      6'b101001 : _zz_shift_i_3_2 = shift_i_map_41;
      6'b101010 : _zz_shift_i_3_2 = shift_i_map_42;
      6'b101011 : _zz_shift_i_3_2 = shift_i_map_43;
      6'b101100 : _zz_shift_i_3_2 = shift_i_map_44;
      6'b101101 : _zz_shift_i_3_2 = shift_i_map_45;
      6'b101110 : _zz_shift_i_3_2 = shift_i_map_46;
      6'b101111 : _zz_shift_i_3_2 = shift_i_map_47;
      6'b110000 : _zz_shift_i_3_2 = shift_i_map_48;
      6'b110001 : _zz_shift_i_3_2 = shift_i_map_49;
      6'b110010 : _zz_shift_i_3_2 = shift_i_map_50;
      6'b110011 : _zz_shift_i_3_2 = shift_i_map_51;
      6'b110100 : _zz_shift_i_3_2 = shift_i_map_52;
      6'b110101 : _zz_shift_i_3_2 = shift_i_map_53;
      6'b110110 : _zz_shift_i_3_2 = shift_i_map_54;
      6'b110111 : _zz_shift_i_3_2 = shift_i_map_55;
      6'b111000 : _zz_shift_i_3_2 = shift_i_map_56;
      6'b111001 : _zz_shift_i_3_2 = shift_i_map_57;
      6'b111010 : _zz_shift_i_3_2 = shift_i_map_58;
      6'b111011 : _zz_shift_i_3_2 = shift_i_map_59;
      6'b111100 : _zz_shift_i_3_2 = shift_i_map_60;
      6'b111101 : _zz_shift_i_3_2 = shift_i_map_61;
      6'b111110 : _zz_shift_i_3_2 = shift_i_map_62;
      default : _zz_shift_i_3_2 = shift_i_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_3_3)
      6'b000000 : _zz_shift_q_3_2 = shift_q_map_0;
      6'b000001 : _zz_shift_q_3_2 = shift_q_map_1;
      6'b000010 : _zz_shift_q_3_2 = shift_q_map_2;
      6'b000011 : _zz_shift_q_3_2 = shift_q_map_3;
      6'b000100 : _zz_shift_q_3_2 = shift_q_map_4;
      6'b000101 : _zz_shift_q_3_2 = shift_q_map_5;
      6'b000110 : _zz_shift_q_3_2 = shift_q_map_6;
      6'b000111 : _zz_shift_q_3_2 = shift_q_map_7;
      6'b001000 : _zz_shift_q_3_2 = shift_q_map_8;
      6'b001001 : _zz_shift_q_3_2 = shift_q_map_9;
      6'b001010 : _zz_shift_q_3_2 = shift_q_map_10;
      6'b001011 : _zz_shift_q_3_2 = shift_q_map_11;
      6'b001100 : _zz_shift_q_3_2 = shift_q_map_12;
      6'b001101 : _zz_shift_q_3_2 = shift_q_map_13;
      6'b001110 : _zz_shift_q_3_2 = shift_q_map_14;
      6'b001111 : _zz_shift_q_3_2 = shift_q_map_15;
      6'b010000 : _zz_shift_q_3_2 = shift_q_map_16;
      6'b010001 : _zz_shift_q_3_2 = shift_q_map_17;
      6'b010010 : _zz_shift_q_3_2 = shift_q_map_18;
      6'b010011 : _zz_shift_q_3_2 = shift_q_map_19;
      6'b010100 : _zz_shift_q_3_2 = shift_q_map_20;
      6'b010101 : _zz_shift_q_3_2 = shift_q_map_21;
      6'b010110 : _zz_shift_q_3_2 = shift_q_map_22;
      6'b010111 : _zz_shift_q_3_2 = shift_q_map_23;
      6'b011000 : _zz_shift_q_3_2 = shift_q_map_24;
      6'b011001 : _zz_shift_q_3_2 = shift_q_map_25;
      6'b011010 : _zz_shift_q_3_2 = shift_q_map_26;
      6'b011011 : _zz_shift_q_3_2 = shift_q_map_27;
      6'b011100 : _zz_shift_q_3_2 = shift_q_map_28;
      6'b011101 : _zz_shift_q_3_2 = shift_q_map_29;
      6'b011110 : _zz_shift_q_3_2 = shift_q_map_30;
      6'b011111 : _zz_shift_q_3_2 = shift_q_map_31;
      6'b100000 : _zz_shift_q_3_2 = shift_q_map_32;
      6'b100001 : _zz_shift_q_3_2 = shift_q_map_33;
      6'b100010 : _zz_shift_q_3_2 = shift_q_map_34;
      6'b100011 : _zz_shift_q_3_2 = shift_q_map_35;
      6'b100100 : _zz_shift_q_3_2 = shift_q_map_36;
      6'b100101 : _zz_shift_q_3_2 = shift_q_map_37;
      6'b100110 : _zz_shift_q_3_2 = shift_q_map_38;
      6'b100111 : _zz_shift_q_3_2 = shift_q_map_39;
      6'b101000 : _zz_shift_q_3_2 = shift_q_map_40;
      6'b101001 : _zz_shift_q_3_2 = shift_q_map_41;
      6'b101010 : _zz_shift_q_3_2 = shift_q_map_42;
      6'b101011 : _zz_shift_q_3_2 = shift_q_map_43;
      6'b101100 : _zz_shift_q_3_2 = shift_q_map_44;
      6'b101101 : _zz_shift_q_3_2 = shift_q_map_45;
      6'b101110 : _zz_shift_q_3_2 = shift_q_map_46;
      6'b101111 : _zz_shift_q_3_2 = shift_q_map_47;
      6'b110000 : _zz_shift_q_3_2 = shift_q_map_48;
      6'b110001 : _zz_shift_q_3_2 = shift_q_map_49;
      6'b110010 : _zz_shift_q_3_2 = shift_q_map_50;
      6'b110011 : _zz_shift_q_3_2 = shift_q_map_51;
      6'b110100 : _zz_shift_q_3_2 = shift_q_map_52;
      6'b110101 : _zz_shift_q_3_2 = shift_q_map_53;
      6'b110110 : _zz_shift_q_3_2 = shift_q_map_54;
      6'b110111 : _zz_shift_q_3_2 = shift_q_map_55;
      6'b111000 : _zz_shift_q_3_2 = shift_q_map_56;
      6'b111001 : _zz_shift_q_3_2 = shift_q_map_57;
      6'b111010 : _zz_shift_q_3_2 = shift_q_map_58;
      6'b111011 : _zz_shift_q_3_2 = shift_q_map_59;
      6'b111100 : _zz_shift_q_3_2 = shift_q_map_60;
      6'b111101 : _zz_shift_q_3_2 = shift_q_map_61;
      6'b111110 : _zz_shift_q_3_2 = shift_q_map_62;
      default : _zz_shift_q_3_2 = shift_q_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_4_3)
      6'b000000 : _zz_shift_i_4_2 = shift_i_map_0;
      6'b000001 : _zz_shift_i_4_2 = shift_i_map_1;
      6'b000010 : _zz_shift_i_4_2 = shift_i_map_2;
      6'b000011 : _zz_shift_i_4_2 = shift_i_map_3;
      6'b000100 : _zz_shift_i_4_2 = shift_i_map_4;
      6'b000101 : _zz_shift_i_4_2 = shift_i_map_5;
      6'b000110 : _zz_shift_i_4_2 = shift_i_map_6;
      6'b000111 : _zz_shift_i_4_2 = shift_i_map_7;
      6'b001000 : _zz_shift_i_4_2 = shift_i_map_8;
      6'b001001 : _zz_shift_i_4_2 = shift_i_map_9;
      6'b001010 : _zz_shift_i_4_2 = shift_i_map_10;
      6'b001011 : _zz_shift_i_4_2 = shift_i_map_11;
      6'b001100 : _zz_shift_i_4_2 = shift_i_map_12;
      6'b001101 : _zz_shift_i_4_2 = shift_i_map_13;
      6'b001110 : _zz_shift_i_4_2 = shift_i_map_14;
      6'b001111 : _zz_shift_i_4_2 = shift_i_map_15;
      6'b010000 : _zz_shift_i_4_2 = shift_i_map_16;
      6'b010001 : _zz_shift_i_4_2 = shift_i_map_17;
      6'b010010 : _zz_shift_i_4_2 = shift_i_map_18;
      6'b010011 : _zz_shift_i_4_2 = shift_i_map_19;
      6'b010100 : _zz_shift_i_4_2 = shift_i_map_20;
      6'b010101 : _zz_shift_i_4_2 = shift_i_map_21;
      6'b010110 : _zz_shift_i_4_2 = shift_i_map_22;
      6'b010111 : _zz_shift_i_4_2 = shift_i_map_23;
      6'b011000 : _zz_shift_i_4_2 = shift_i_map_24;
      6'b011001 : _zz_shift_i_4_2 = shift_i_map_25;
      6'b011010 : _zz_shift_i_4_2 = shift_i_map_26;
      6'b011011 : _zz_shift_i_4_2 = shift_i_map_27;
      6'b011100 : _zz_shift_i_4_2 = shift_i_map_28;
      6'b011101 : _zz_shift_i_4_2 = shift_i_map_29;
      6'b011110 : _zz_shift_i_4_2 = shift_i_map_30;
      6'b011111 : _zz_shift_i_4_2 = shift_i_map_31;
      6'b100000 : _zz_shift_i_4_2 = shift_i_map_32;
      6'b100001 : _zz_shift_i_4_2 = shift_i_map_33;
      6'b100010 : _zz_shift_i_4_2 = shift_i_map_34;
      6'b100011 : _zz_shift_i_4_2 = shift_i_map_35;
      6'b100100 : _zz_shift_i_4_2 = shift_i_map_36;
      6'b100101 : _zz_shift_i_4_2 = shift_i_map_37;
      6'b100110 : _zz_shift_i_4_2 = shift_i_map_38;
      6'b100111 : _zz_shift_i_4_2 = shift_i_map_39;
      6'b101000 : _zz_shift_i_4_2 = shift_i_map_40;
      6'b101001 : _zz_shift_i_4_2 = shift_i_map_41;
      6'b101010 : _zz_shift_i_4_2 = shift_i_map_42;
      6'b101011 : _zz_shift_i_4_2 = shift_i_map_43;
      6'b101100 : _zz_shift_i_4_2 = shift_i_map_44;
      6'b101101 : _zz_shift_i_4_2 = shift_i_map_45;
      6'b101110 : _zz_shift_i_4_2 = shift_i_map_46;
      6'b101111 : _zz_shift_i_4_2 = shift_i_map_47;
      6'b110000 : _zz_shift_i_4_2 = shift_i_map_48;
      6'b110001 : _zz_shift_i_4_2 = shift_i_map_49;
      6'b110010 : _zz_shift_i_4_2 = shift_i_map_50;
      6'b110011 : _zz_shift_i_4_2 = shift_i_map_51;
      6'b110100 : _zz_shift_i_4_2 = shift_i_map_52;
      6'b110101 : _zz_shift_i_4_2 = shift_i_map_53;
      6'b110110 : _zz_shift_i_4_2 = shift_i_map_54;
      6'b110111 : _zz_shift_i_4_2 = shift_i_map_55;
      6'b111000 : _zz_shift_i_4_2 = shift_i_map_56;
      6'b111001 : _zz_shift_i_4_2 = shift_i_map_57;
      6'b111010 : _zz_shift_i_4_2 = shift_i_map_58;
      6'b111011 : _zz_shift_i_4_2 = shift_i_map_59;
      6'b111100 : _zz_shift_i_4_2 = shift_i_map_60;
      6'b111101 : _zz_shift_i_4_2 = shift_i_map_61;
      6'b111110 : _zz_shift_i_4_2 = shift_i_map_62;
      default : _zz_shift_i_4_2 = shift_i_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_4_3)
      6'b000000 : _zz_shift_q_4_2 = shift_q_map_0;
      6'b000001 : _zz_shift_q_4_2 = shift_q_map_1;
      6'b000010 : _zz_shift_q_4_2 = shift_q_map_2;
      6'b000011 : _zz_shift_q_4_2 = shift_q_map_3;
      6'b000100 : _zz_shift_q_4_2 = shift_q_map_4;
      6'b000101 : _zz_shift_q_4_2 = shift_q_map_5;
      6'b000110 : _zz_shift_q_4_2 = shift_q_map_6;
      6'b000111 : _zz_shift_q_4_2 = shift_q_map_7;
      6'b001000 : _zz_shift_q_4_2 = shift_q_map_8;
      6'b001001 : _zz_shift_q_4_2 = shift_q_map_9;
      6'b001010 : _zz_shift_q_4_2 = shift_q_map_10;
      6'b001011 : _zz_shift_q_4_2 = shift_q_map_11;
      6'b001100 : _zz_shift_q_4_2 = shift_q_map_12;
      6'b001101 : _zz_shift_q_4_2 = shift_q_map_13;
      6'b001110 : _zz_shift_q_4_2 = shift_q_map_14;
      6'b001111 : _zz_shift_q_4_2 = shift_q_map_15;
      6'b010000 : _zz_shift_q_4_2 = shift_q_map_16;
      6'b010001 : _zz_shift_q_4_2 = shift_q_map_17;
      6'b010010 : _zz_shift_q_4_2 = shift_q_map_18;
      6'b010011 : _zz_shift_q_4_2 = shift_q_map_19;
      6'b010100 : _zz_shift_q_4_2 = shift_q_map_20;
      6'b010101 : _zz_shift_q_4_2 = shift_q_map_21;
      6'b010110 : _zz_shift_q_4_2 = shift_q_map_22;
      6'b010111 : _zz_shift_q_4_2 = shift_q_map_23;
      6'b011000 : _zz_shift_q_4_2 = shift_q_map_24;
      6'b011001 : _zz_shift_q_4_2 = shift_q_map_25;
      6'b011010 : _zz_shift_q_4_2 = shift_q_map_26;
      6'b011011 : _zz_shift_q_4_2 = shift_q_map_27;
      6'b011100 : _zz_shift_q_4_2 = shift_q_map_28;
      6'b011101 : _zz_shift_q_4_2 = shift_q_map_29;
      6'b011110 : _zz_shift_q_4_2 = shift_q_map_30;
      6'b011111 : _zz_shift_q_4_2 = shift_q_map_31;
      6'b100000 : _zz_shift_q_4_2 = shift_q_map_32;
      6'b100001 : _zz_shift_q_4_2 = shift_q_map_33;
      6'b100010 : _zz_shift_q_4_2 = shift_q_map_34;
      6'b100011 : _zz_shift_q_4_2 = shift_q_map_35;
      6'b100100 : _zz_shift_q_4_2 = shift_q_map_36;
      6'b100101 : _zz_shift_q_4_2 = shift_q_map_37;
      6'b100110 : _zz_shift_q_4_2 = shift_q_map_38;
      6'b100111 : _zz_shift_q_4_2 = shift_q_map_39;
      6'b101000 : _zz_shift_q_4_2 = shift_q_map_40;
      6'b101001 : _zz_shift_q_4_2 = shift_q_map_41;
      6'b101010 : _zz_shift_q_4_2 = shift_q_map_42;
      6'b101011 : _zz_shift_q_4_2 = shift_q_map_43;
      6'b101100 : _zz_shift_q_4_2 = shift_q_map_44;
      6'b101101 : _zz_shift_q_4_2 = shift_q_map_45;
      6'b101110 : _zz_shift_q_4_2 = shift_q_map_46;
      6'b101111 : _zz_shift_q_4_2 = shift_q_map_47;
      6'b110000 : _zz_shift_q_4_2 = shift_q_map_48;
      6'b110001 : _zz_shift_q_4_2 = shift_q_map_49;
      6'b110010 : _zz_shift_q_4_2 = shift_q_map_50;
      6'b110011 : _zz_shift_q_4_2 = shift_q_map_51;
      6'b110100 : _zz_shift_q_4_2 = shift_q_map_52;
      6'b110101 : _zz_shift_q_4_2 = shift_q_map_53;
      6'b110110 : _zz_shift_q_4_2 = shift_q_map_54;
      6'b110111 : _zz_shift_q_4_2 = shift_q_map_55;
      6'b111000 : _zz_shift_q_4_2 = shift_q_map_56;
      6'b111001 : _zz_shift_q_4_2 = shift_q_map_57;
      6'b111010 : _zz_shift_q_4_2 = shift_q_map_58;
      6'b111011 : _zz_shift_q_4_2 = shift_q_map_59;
      6'b111100 : _zz_shift_q_4_2 = shift_q_map_60;
      6'b111101 : _zz_shift_q_4_2 = shift_q_map_61;
      6'b111110 : _zz_shift_q_4_2 = shift_q_map_62;
      default : _zz_shift_q_4_2 = shift_q_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_5_3)
      6'b000000 : _zz_shift_i_5_2 = shift_i_map_0;
      6'b000001 : _zz_shift_i_5_2 = shift_i_map_1;
      6'b000010 : _zz_shift_i_5_2 = shift_i_map_2;
      6'b000011 : _zz_shift_i_5_2 = shift_i_map_3;
      6'b000100 : _zz_shift_i_5_2 = shift_i_map_4;
      6'b000101 : _zz_shift_i_5_2 = shift_i_map_5;
      6'b000110 : _zz_shift_i_5_2 = shift_i_map_6;
      6'b000111 : _zz_shift_i_5_2 = shift_i_map_7;
      6'b001000 : _zz_shift_i_5_2 = shift_i_map_8;
      6'b001001 : _zz_shift_i_5_2 = shift_i_map_9;
      6'b001010 : _zz_shift_i_5_2 = shift_i_map_10;
      6'b001011 : _zz_shift_i_5_2 = shift_i_map_11;
      6'b001100 : _zz_shift_i_5_2 = shift_i_map_12;
      6'b001101 : _zz_shift_i_5_2 = shift_i_map_13;
      6'b001110 : _zz_shift_i_5_2 = shift_i_map_14;
      6'b001111 : _zz_shift_i_5_2 = shift_i_map_15;
      6'b010000 : _zz_shift_i_5_2 = shift_i_map_16;
      6'b010001 : _zz_shift_i_5_2 = shift_i_map_17;
      6'b010010 : _zz_shift_i_5_2 = shift_i_map_18;
      6'b010011 : _zz_shift_i_5_2 = shift_i_map_19;
      6'b010100 : _zz_shift_i_5_2 = shift_i_map_20;
      6'b010101 : _zz_shift_i_5_2 = shift_i_map_21;
      6'b010110 : _zz_shift_i_5_2 = shift_i_map_22;
      6'b010111 : _zz_shift_i_5_2 = shift_i_map_23;
      6'b011000 : _zz_shift_i_5_2 = shift_i_map_24;
      6'b011001 : _zz_shift_i_5_2 = shift_i_map_25;
      6'b011010 : _zz_shift_i_5_2 = shift_i_map_26;
      6'b011011 : _zz_shift_i_5_2 = shift_i_map_27;
      6'b011100 : _zz_shift_i_5_2 = shift_i_map_28;
      6'b011101 : _zz_shift_i_5_2 = shift_i_map_29;
      6'b011110 : _zz_shift_i_5_2 = shift_i_map_30;
      6'b011111 : _zz_shift_i_5_2 = shift_i_map_31;
      6'b100000 : _zz_shift_i_5_2 = shift_i_map_32;
      6'b100001 : _zz_shift_i_5_2 = shift_i_map_33;
      6'b100010 : _zz_shift_i_5_2 = shift_i_map_34;
      6'b100011 : _zz_shift_i_5_2 = shift_i_map_35;
      6'b100100 : _zz_shift_i_5_2 = shift_i_map_36;
      6'b100101 : _zz_shift_i_5_2 = shift_i_map_37;
      6'b100110 : _zz_shift_i_5_2 = shift_i_map_38;
      6'b100111 : _zz_shift_i_5_2 = shift_i_map_39;
      6'b101000 : _zz_shift_i_5_2 = shift_i_map_40;
      6'b101001 : _zz_shift_i_5_2 = shift_i_map_41;
      6'b101010 : _zz_shift_i_5_2 = shift_i_map_42;
      6'b101011 : _zz_shift_i_5_2 = shift_i_map_43;
      6'b101100 : _zz_shift_i_5_2 = shift_i_map_44;
      6'b101101 : _zz_shift_i_5_2 = shift_i_map_45;
      6'b101110 : _zz_shift_i_5_2 = shift_i_map_46;
      6'b101111 : _zz_shift_i_5_2 = shift_i_map_47;
      6'b110000 : _zz_shift_i_5_2 = shift_i_map_48;
      6'b110001 : _zz_shift_i_5_2 = shift_i_map_49;
      6'b110010 : _zz_shift_i_5_2 = shift_i_map_50;
      6'b110011 : _zz_shift_i_5_2 = shift_i_map_51;
      6'b110100 : _zz_shift_i_5_2 = shift_i_map_52;
      6'b110101 : _zz_shift_i_5_2 = shift_i_map_53;
      6'b110110 : _zz_shift_i_5_2 = shift_i_map_54;
      6'b110111 : _zz_shift_i_5_2 = shift_i_map_55;
      6'b111000 : _zz_shift_i_5_2 = shift_i_map_56;
      6'b111001 : _zz_shift_i_5_2 = shift_i_map_57;
      6'b111010 : _zz_shift_i_5_2 = shift_i_map_58;
      6'b111011 : _zz_shift_i_5_2 = shift_i_map_59;
      6'b111100 : _zz_shift_i_5_2 = shift_i_map_60;
      6'b111101 : _zz_shift_i_5_2 = shift_i_map_61;
      6'b111110 : _zz_shift_i_5_2 = shift_i_map_62;
      default : _zz_shift_i_5_2 = shift_i_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_5_3)
      6'b000000 : _zz_shift_q_5_2 = shift_q_map_0;
      6'b000001 : _zz_shift_q_5_2 = shift_q_map_1;
      6'b000010 : _zz_shift_q_5_2 = shift_q_map_2;
      6'b000011 : _zz_shift_q_5_2 = shift_q_map_3;
      6'b000100 : _zz_shift_q_5_2 = shift_q_map_4;
      6'b000101 : _zz_shift_q_5_2 = shift_q_map_5;
      6'b000110 : _zz_shift_q_5_2 = shift_q_map_6;
      6'b000111 : _zz_shift_q_5_2 = shift_q_map_7;
      6'b001000 : _zz_shift_q_5_2 = shift_q_map_8;
      6'b001001 : _zz_shift_q_5_2 = shift_q_map_9;
      6'b001010 : _zz_shift_q_5_2 = shift_q_map_10;
      6'b001011 : _zz_shift_q_5_2 = shift_q_map_11;
      6'b001100 : _zz_shift_q_5_2 = shift_q_map_12;
      6'b001101 : _zz_shift_q_5_2 = shift_q_map_13;
      6'b001110 : _zz_shift_q_5_2 = shift_q_map_14;
      6'b001111 : _zz_shift_q_5_2 = shift_q_map_15;
      6'b010000 : _zz_shift_q_5_2 = shift_q_map_16;
      6'b010001 : _zz_shift_q_5_2 = shift_q_map_17;
      6'b010010 : _zz_shift_q_5_2 = shift_q_map_18;
      6'b010011 : _zz_shift_q_5_2 = shift_q_map_19;
      6'b010100 : _zz_shift_q_5_2 = shift_q_map_20;
      6'b010101 : _zz_shift_q_5_2 = shift_q_map_21;
      6'b010110 : _zz_shift_q_5_2 = shift_q_map_22;
      6'b010111 : _zz_shift_q_5_2 = shift_q_map_23;
      6'b011000 : _zz_shift_q_5_2 = shift_q_map_24;
      6'b011001 : _zz_shift_q_5_2 = shift_q_map_25;
      6'b011010 : _zz_shift_q_5_2 = shift_q_map_26;
      6'b011011 : _zz_shift_q_5_2 = shift_q_map_27;
      6'b011100 : _zz_shift_q_5_2 = shift_q_map_28;
      6'b011101 : _zz_shift_q_5_2 = shift_q_map_29;
      6'b011110 : _zz_shift_q_5_2 = shift_q_map_30;
      6'b011111 : _zz_shift_q_5_2 = shift_q_map_31;
      6'b100000 : _zz_shift_q_5_2 = shift_q_map_32;
      6'b100001 : _zz_shift_q_5_2 = shift_q_map_33;
      6'b100010 : _zz_shift_q_5_2 = shift_q_map_34;
      6'b100011 : _zz_shift_q_5_2 = shift_q_map_35;
      6'b100100 : _zz_shift_q_5_2 = shift_q_map_36;
      6'b100101 : _zz_shift_q_5_2 = shift_q_map_37;
      6'b100110 : _zz_shift_q_5_2 = shift_q_map_38;
      6'b100111 : _zz_shift_q_5_2 = shift_q_map_39;
      6'b101000 : _zz_shift_q_5_2 = shift_q_map_40;
      6'b101001 : _zz_shift_q_5_2 = shift_q_map_41;
      6'b101010 : _zz_shift_q_5_2 = shift_q_map_42;
      6'b101011 : _zz_shift_q_5_2 = shift_q_map_43;
      6'b101100 : _zz_shift_q_5_2 = shift_q_map_44;
      6'b101101 : _zz_shift_q_5_2 = shift_q_map_45;
      6'b101110 : _zz_shift_q_5_2 = shift_q_map_46;
      6'b101111 : _zz_shift_q_5_2 = shift_q_map_47;
      6'b110000 : _zz_shift_q_5_2 = shift_q_map_48;
      6'b110001 : _zz_shift_q_5_2 = shift_q_map_49;
      6'b110010 : _zz_shift_q_5_2 = shift_q_map_50;
      6'b110011 : _zz_shift_q_5_2 = shift_q_map_51;
      6'b110100 : _zz_shift_q_5_2 = shift_q_map_52;
      6'b110101 : _zz_shift_q_5_2 = shift_q_map_53;
      6'b110110 : _zz_shift_q_5_2 = shift_q_map_54;
      6'b110111 : _zz_shift_q_5_2 = shift_q_map_55;
      6'b111000 : _zz_shift_q_5_2 = shift_q_map_56;
      6'b111001 : _zz_shift_q_5_2 = shift_q_map_57;
      6'b111010 : _zz_shift_q_5_2 = shift_q_map_58;
      6'b111011 : _zz_shift_q_5_2 = shift_q_map_59;
      6'b111100 : _zz_shift_q_5_2 = shift_q_map_60;
      6'b111101 : _zz_shift_q_5_2 = shift_q_map_61;
      6'b111110 : _zz_shift_q_5_2 = shift_q_map_62;
      default : _zz_shift_q_5_2 = shift_q_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_6_3)
      6'b000000 : _zz_shift_i_6_2 = shift_i_map_0;
      6'b000001 : _zz_shift_i_6_2 = shift_i_map_1;
      6'b000010 : _zz_shift_i_6_2 = shift_i_map_2;
      6'b000011 : _zz_shift_i_6_2 = shift_i_map_3;
      6'b000100 : _zz_shift_i_6_2 = shift_i_map_4;
      6'b000101 : _zz_shift_i_6_2 = shift_i_map_5;
      6'b000110 : _zz_shift_i_6_2 = shift_i_map_6;
      6'b000111 : _zz_shift_i_6_2 = shift_i_map_7;
      6'b001000 : _zz_shift_i_6_2 = shift_i_map_8;
      6'b001001 : _zz_shift_i_6_2 = shift_i_map_9;
      6'b001010 : _zz_shift_i_6_2 = shift_i_map_10;
      6'b001011 : _zz_shift_i_6_2 = shift_i_map_11;
      6'b001100 : _zz_shift_i_6_2 = shift_i_map_12;
      6'b001101 : _zz_shift_i_6_2 = shift_i_map_13;
      6'b001110 : _zz_shift_i_6_2 = shift_i_map_14;
      6'b001111 : _zz_shift_i_6_2 = shift_i_map_15;
      6'b010000 : _zz_shift_i_6_2 = shift_i_map_16;
      6'b010001 : _zz_shift_i_6_2 = shift_i_map_17;
      6'b010010 : _zz_shift_i_6_2 = shift_i_map_18;
      6'b010011 : _zz_shift_i_6_2 = shift_i_map_19;
      6'b010100 : _zz_shift_i_6_2 = shift_i_map_20;
      6'b010101 : _zz_shift_i_6_2 = shift_i_map_21;
      6'b010110 : _zz_shift_i_6_2 = shift_i_map_22;
      6'b010111 : _zz_shift_i_6_2 = shift_i_map_23;
      6'b011000 : _zz_shift_i_6_2 = shift_i_map_24;
      6'b011001 : _zz_shift_i_6_2 = shift_i_map_25;
      6'b011010 : _zz_shift_i_6_2 = shift_i_map_26;
      6'b011011 : _zz_shift_i_6_2 = shift_i_map_27;
      6'b011100 : _zz_shift_i_6_2 = shift_i_map_28;
      6'b011101 : _zz_shift_i_6_2 = shift_i_map_29;
      6'b011110 : _zz_shift_i_6_2 = shift_i_map_30;
      6'b011111 : _zz_shift_i_6_2 = shift_i_map_31;
      6'b100000 : _zz_shift_i_6_2 = shift_i_map_32;
      6'b100001 : _zz_shift_i_6_2 = shift_i_map_33;
      6'b100010 : _zz_shift_i_6_2 = shift_i_map_34;
      6'b100011 : _zz_shift_i_6_2 = shift_i_map_35;
      6'b100100 : _zz_shift_i_6_2 = shift_i_map_36;
      6'b100101 : _zz_shift_i_6_2 = shift_i_map_37;
      6'b100110 : _zz_shift_i_6_2 = shift_i_map_38;
      6'b100111 : _zz_shift_i_6_2 = shift_i_map_39;
      6'b101000 : _zz_shift_i_6_2 = shift_i_map_40;
      6'b101001 : _zz_shift_i_6_2 = shift_i_map_41;
      6'b101010 : _zz_shift_i_6_2 = shift_i_map_42;
      6'b101011 : _zz_shift_i_6_2 = shift_i_map_43;
      6'b101100 : _zz_shift_i_6_2 = shift_i_map_44;
      6'b101101 : _zz_shift_i_6_2 = shift_i_map_45;
      6'b101110 : _zz_shift_i_6_2 = shift_i_map_46;
      6'b101111 : _zz_shift_i_6_2 = shift_i_map_47;
      6'b110000 : _zz_shift_i_6_2 = shift_i_map_48;
      6'b110001 : _zz_shift_i_6_2 = shift_i_map_49;
      6'b110010 : _zz_shift_i_6_2 = shift_i_map_50;
      6'b110011 : _zz_shift_i_6_2 = shift_i_map_51;
      6'b110100 : _zz_shift_i_6_2 = shift_i_map_52;
      6'b110101 : _zz_shift_i_6_2 = shift_i_map_53;
      6'b110110 : _zz_shift_i_6_2 = shift_i_map_54;
      6'b110111 : _zz_shift_i_6_2 = shift_i_map_55;
      6'b111000 : _zz_shift_i_6_2 = shift_i_map_56;
      6'b111001 : _zz_shift_i_6_2 = shift_i_map_57;
      6'b111010 : _zz_shift_i_6_2 = shift_i_map_58;
      6'b111011 : _zz_shift_i_6_2 = shift_i_map_59;
      6'b111100 : _zz_shift_i_6_2 = shift_i_map_60;
      6'b111101 : _zz_shift_i_6_2 = shift_i_map_61;
      6'b111110 : _zz_shift_i_6_2 = shift_i_map_62;
      default : _zz_shift_i_6_2 = shift_i_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_6_3)
      6'b000000 : _zz_shift_q_6_2 = shift_q_map_0;
      6'b000001 : _zz_shift_q_6_2 = shift_q_map_1;
      6'b000010 : _zz_shift_q_6_2 = shift_q_map_2;
      6'b000011 : _zz_shift_q_6_2 = shift_q_map_3;
      6'b000100 : _zz_shift_q_6_2 = shift_q_map_4;
      6'b000101 : _zz_shift_q_6_2 = shift_q_map_5;
      6'b000110 : _zz_shift_q_6_2 = shift_q_map_6;
      6'b000111 : _zz_shift_q_6_2 = shift_q_map_7;
      6'b001000 : _zz_shift_q_6_2 = shift_q_map_8;
      6'b001001 : _zz_shift_q_6_2 = shift_q_map_9;
      6'b001010 : _zz_shift_q_6_2 = shift_q_map_10;
      6'b001011 : _zz_shift_q_6_2 = shift_q_map_11;
      6'b001100 : _zz_shift_q_6_2 = shift_q_map_12;
      6'b001101 : _zz_shift_q_6_2 = shift_q_map_13;
      6'b001110 : _zz_shift_q_6_2 = shift_q_map_14;
      6'b001111 : _zz_shift_q_6_2 = shift_q_map_15;
      6'b010000 : _zz_shift_q_6_2 = shift_q_map_16;
      6'b010001 : _zz_shift_q_6_2 = shift_q_map_17;
      6'b010010 : _zz_shift_q_6_2 = shift_q_map_18;
      6'b010011 : _zz_shift_q_6_2 = shift_q_map_19;
      6'b010100 : _zz_shift_q_6_2 = shift_q_map_20;
      6'b010101 : _zz_shift_q_6_2 = shift_q_map_21;
      6'b010110 : _zz_shift_q_6_2 = shift_q_map_22;
      6'b010111 : _zz_shift_q_6_2 = shift_q_map_23;
      6'b011000 : _zz_shift_q_6_2 = shift_q_map_24;
      6'b011001 : _zz_shift_q_6_2 = shift_q_map_25;
      6'b011010 : _zz_shift_q_6_2 = shift_q_map_26;
      6'b011011 : _zz_shift_q_6_2 = shift_q_map_27;
      6'b011100 : _zz_shift_q_6_2 = shift_q_map_28;
      6'b011101 : _zz_shift_q_6_2 = shift_q_map_29;
      6'b011110 : _zz_shift_q_6_2 = shift_q_map_30;
      6'b011111 : _zz_shift_q_6_2 = shift_q_map_31;
      6'b100000 : _zz_shift_q_6_2 = shift_q_map_32;
      6'b100001 : _zz_shift_q_6_2 = shift_q_map_33;
      6'b100010 : _zz_shift_q_6_2 = shift_q_map_34;
      6'b100011 : _zz_shift_q_6_2 = shift_q_map_35;
      6'b100100 : _zz_shift_q_6_2 = shift_q_map_36;
      6'b100101 : _zz_shift_q_6_2 = shift_q_map_37;
      6'b100110 : _zz_shift_q_6_2 = shift_q_map_38;
      6'b100111 : _zz_shift_q_6_2 = shift_q_map_39;
      6'b101000 : _zz_shift_q_6_2 = shift_q_map_40;
      6'b101001 : _zz_shift_q_6_2 = shift_q_map_41;
      6'b101010 : _zz_shift_q_6_2 = shift_q_map_42;
      6'b101011 : _zz_shift_q_6_2 = shift_q_map_43;
      6'b101100 : _zz_shift_q_6_2 = shift_q_map_44;
      6'b101101 : _zz_shift_q_6_2 = shift_q_map_45;
      6'b101110 : _zz_shift_q_6_2 = shift_q_map_46;
      6'b101111 : _zz_shift_q_6_2 = shift_q_map_47;
      6'b110000 : _zz_shift_q_6_2 = shift_q_map_48;
      6'b110001 : _zz_shift_q_6_2 = shift_q_map_49;
      6'b110010 : _zz_shift_q_6_2 = shift_q_map_50;
      6'b110011 : _zz_shift_q_6_2 = shift_q_map_51;
      6'b110100 : _zz_shift_q_6_2 = shift_q_map_52;
      6'b110101 : _zz_shift_q_6_2 = shift_q_map_53;
      6'b110110 : _zz_shift_q_6_2 = shift_q_map_54;
      6'b110111 : _zz_shift_q_6_2 = shift_q_map_55;
      6'b111000 : _zz_shift_q_6_2 = shift_q_map_56;
      6'b111001 : _zz_shift_q_6_2 = shift_q_map_57;
      6'b111010 : _zz_shift_q_6_2 = shift_q_map_58;
      6'b111011 : _zz_shift_q_6_2 = shift_q_map_59;
      6'b111100 : _zz_shift_q_6_2 = shift_q_map_60;
      6'b111101 : _zz_shift_q_6_2 = shift_q_map_61;
      6'b111110 : _zz_shift_q_6_2 = shift_q_map_62;
      default : _zz_shift_q_6_2 = shift_q_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_7_3)
      6'b000000 : _zz_shift_i_7_2 = shift_i_map_0;
      6'b000001 : _zz_shift_i_7_2 = shift_i_map_1;
      6'b000010 : _zz_shift_i_7_2 = shift_i_map_2;
      6'b000011 : _zz_shift_i_7_2 = shift_i_map_3;
      6'b000100 : _zz_shift_i_7_2 = shift_i_map_4;
      6'b000101 : _zz_shift_i_7_2 = shift_i_map_5;
      6'b000110 : _zz_shift_i_7_2 = shift_i_map_6;
      6'b000111 : _zz_shift_i_7_2 = shift_i_map_7;
      6'b001000 : _zz_shift_i_7_2 = shift_i_map_8;
      6'b001001 : _zz_shift_i_7_2 = shift_i_map_9;
      6'b001010 : _zz_shift_i_7_2 = shift_i_map_10;
      6'b001011 : _zz_shift_i_7_2 = shift_i_map_11;
      6'b001100 : _zz_shift_i_7_2 = shift_i_map_12;
      6'b001101 : _zz_shift_i_7_2 = shift_i_map_13;
      6'b001110 : _zz_shift_i_7_2 = shift_i_map_14;
      6'b001111 : _zz_shift_i_7_2 = shift_i_map_15;
      6'b010000 : _zz_shift_i_7_2 = shift_i_map_16;
      6'b010001 : _zz_shift_i_7_2 = shift_i_map_17;
      6'b010010 : _zz_shift_i_7_2 = shift_i_map_18;
      6'b010011 : _zz_shift_i_7_2 = shift_i_map_19;
      6'b010100 : _zz_shift_i_7_2 = shift_i_map_20;
      6'b010101 : _zz_shift_i_7_2 = shift_i_map_21;
      6'b010110 : _zz_shift_i_7_2 = shift_i_map_22;
      6'b010111 : _zz_shift_i_7_2 = shift_i_map_23;
      6'b011000 : _zz_shift_i_7_2 = shift_i_map_24;
      6'b011001 : _zz_shift_i_7_2 = shift_i_map_25;
      6'b011010 : _zz_shift_i_7_2 = shift_i_map_26;
      6'b011011 : _zz_shift_i_7_2 = shift_i_map_27;
      6'b011100 : _zz_shift_i_7_2 = shift_i_map_28;
      6'b011101 : _zz_shift_i_7_2 = shift_i_map_29;
      6'b011110 : _zz_shift_i_7_2 = shift_i_map_30;
      6'b011111 : _zz_shift_i_7_2 = shift_i_map_31;
      6'b100000 : _zz_shift_i_7_2 = shift_i_map_32;
      6'b100001 : _zz_shift_i_7_2 = shift_i_map_33;
      6'b100010 : _zz_shift_i_7_2 = shift_i_map_34;
      6'b100011 : _zz_shift_i_7_2 = shift_i_map_35;
      6'b100100 : _zz_shift_i_7_2 = shift_i_map_36;
      6'b100101 : _zz_shift_i_7_2 = shift_i_map_37;
      6'b100110 : _zz_shift_i_7_2 = shift_i_map_38;
      6'b100111 : _zz_shift_i_7_2 = shift_i_map_39;
      6'b101000 : _zz_shift_i_7_2 = shift_i_map_40;
      6'b101001 : _zz_shift_i_7_2 = shift_i_map_41;
      6'b101010 : _zz_shift_i_7_2 = shift_i_map_42;
      6'b101011 : _zz_shift_i_7_2 = shift_i_map_43;
      6'b101100 : _zz_shift_i_7_2 = shift_i_map_44;
      6'b101101 : _zz_shift_i_7_2 = shift_i_map_45;
      6'b101110 : _zz_shift_i_7_2 = shift_i_map_46;
      6'b101111 : _zz_shift_i_7_2 = shift_i_map_47;
      6'b110000 : _zz_shift_i_7_2 = shift_i_map_48;
      6'b110001 : _zz_shift_i_7_2 = shift_i_map_49;
      6'b110010 : _zz_shift_i_7_2 = shift_i_map_50;
      6'b110011 : _zz_shift_i_7_2 = shift_i_map_51;
      6'b110100 : _zz_shift_i_7_2 = shift_i_map_52;
      6'b110101 : _zz_shift_i_7_2 = shift_i_map_53;
      6'b110110 : _zz_shift_i_7_2 = shift_i_map_54;
      6'b110111 : _zz_shift_i_7_2 = shift_i_map_55;
      6'b111000 : _zz_shift_i_7_2 = shift_i_map_56;
      6'b111001 : _zz_shift_i_7_2 = shift_i_map_57;
      6'b111010 : _zz_shift_i_7_2 = shift_i_map_58;
      6'b111011 : _zz_shift_i_7_2 = shift_i_map_59;
      6'b111100 : _zz_shift_i_7_2 = shift_i_map_60;
      6'b111101 : _zz_shift_i_7_2 = shift_i_map_61;
      6'b111110 : _zz_shift_i_7_2 = shift_i_map_62;
      default : _zz_shift_i_7_2 = shift_i_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_7_3)
      6'b000000 : _zz_shift_q_7_2 = shift_q_map_0;
      6'b000001 : _zz_shift_q_7_2 = shift_q_map_1;
      6'b000010 : _zz_shift_q_7_2 = shift_q_map_2;
      6'b000011 : _zz_shift_q_7_2 = shift_q_map_3;
      6'b000100 : _zz_shift_q_7_2 = shift_q_map_4;
      6'b000101 : _zz_shift_q_7_2 = shift_q_map_5;
      6'b000110 : _zz_shift_q_7_2 = shift_q_map_6;
      6'b000111 : _zz_shift_q_7_2 = shift_q_map_7;
      6'b001000 : _zz_shift_q_7_2 = shift_q_map_8;
      6'b001001 : _zz_shift_q_7_2 = shift_q_map_9;
      6'b001010 : _zz_shift_q_7_2 = shift_q_map_10;
      6'b001011 : _zz_shift_q_7_2 = shift_q_map_11;
      6'b001100 : _zz_shift_q_7_2 = shift_q_map_12;
      6'b001101 : _zz_shift_q_7_2 = shift_q_map_13;
      6'b001110 : _zz_shift_q_7_2 = shift_q_map_14;
      6'b001111 : _zz_shift_q_7_2 = shift_q_map_15;
      6'b010000 : _zz_shift_q_7_2 = shift_q_map_16;
      6'b010001 : _zz_shift_q_7_2 = shift_q_map_17;
      6'b010010 : _zz_shift_q_7_2 = shift_q_map_18;
      6'b010011 : _zz_shift_q_7_2 = shift_q_map_19;
      6'b010100 : _zz_shift_q_7_2 = shift_q_map_20;
      6'b010101 : _zz_shift_q_7_2 = shift_q_map_21;
      6'b010110 : _zz_shift_q_7_2 = shift_q_map_22;
      6'b010111 : _zz_shift_q_7_2 = shift_q_map_23;
      6'b011000 : _zz_shift_q_7_2 = shift_q_map_24;
      6'b011001 : _zz_shift_q_7_2 = shift_q_map_25;
      6'b011010 : _zz_shift_q_7_2 = shift_q_map_26;
      6'b011011 : _zz_shift_q_7_2 = shift_q_map_27;
      6'b011100 : _zz_shift_q_7_2 = shift_q_map_28;
      6'b011101 : _zz_shift_q_7_2 = shift_q_map_29;
      6'b011110 : _zz_shift_q_7_2 = shift_q_map_30;
      6'b011111 : _zz_shift_q_7_2 = shift_q_map_31;
      6'b100000 : _zz_shift_q_7_2 = shift_q_map_32;
      6'b100001 : _zz_shift_q_7_2 = shift_q_map_33;
      6'b100010 : _zz_shift_q_7_2 = shift_q_map_34;
      6'b100011 : _zz_shift_q_7_2 = shift_q_map_35;
      6'b100100 : _zz_shift_q_7_2 = shift_q_map_36;
      6'b100101 : _zz_shift_q_7_2 = shift_q_map_37;
      6'b100110 : _zz_shift_q_7_2 = shift_q_map_38;
      6'b100111 : _zz_shift_q_7_2 = shift_q_map_39;
      6'b101000 : _zz_shift_q_7_2 = shift_q_map_40;
      6'b101001 : _zz_shift_q_7_2 = shift_q_map_41;
      6'b101010 : _zz_shift_q_7_2 = shift_q_map_42;
      6'b101011 : _zz_shift_q_7_2 = shift_q_map_43;
      6'b101100 : _zz_shift_q_7_2 = shift_q_map_44;
      6'b101101 : _zz_shift_q_7_2 = shift_q_map_45;
      6'b101110 : _zz_shift_q_7_2 = shift_q_map_46;
      6'b101111 : _zz_shift_q_7_2 = shift_q_map_47;
      6'b110000 : _zz_shift_q_7_2 = shift_q_map_48;
      6'b110001 : _zz_shift_q_7_2 = shift_q_map_49;
      6'b110010 : _zz_shift_q_7_2 = shift_q_map_50;
      6'b110011 : _zz_shift_q_7_2 = shift_q_map_51;
      6'b110100 : _zz_shift_q_7_2 = shift_q_map_52;
      6'b110101 : _zz_shift_q_7_2 = shift_q_map_53;
      6'b110110 : _zz_shift_q_7_2 = shift_q_map_54;
      6'b110111 : _zz_shift_q_7_2 = shift_q_map_55;
      6'b111000 : _zz_shift_q_7_2 = shift_q_map_56;
      6'b111001 : _zz_shift_q_7_2 = shift_q_map_57;
      6'b111010 : _zz_shift_q_7_2 = shift_q_map_58;
      6'b111011 : _zz_shift_q_7_2 = shift_q_map_59;
      6'b111100 : _zz_shift_q_7_2 = shift_q_map_60;
      6'b111101 : _zz_shift_q_7_2 = shift_q_map_61;
      6'b111110 : _zz_shift_q_7_2 = shift_q_map_62;
      default : _zz_shift_q_7_2 = shift_q_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_0_5)
      6'b000000 : _zz_shift_i_0_4 = shift_i_map_0;
      6'b000001 : _zz_shift_i_0_4 = shift_i_map_1;
      6'b000010 : _zz_shift_i_0_4 = shift_i_map_2;
      6'b000011 : _zz_shift_i_0_4 = shift_i_map_3;
      6'b000100 : _zz_shift_i_0_4 = shift_i_map_4;
      6'b000101 : _zz_shift_i_0_4 = shift_i_map_5;
      6'b000110 : _zz_shift_i_0_4 = shift_i_map_6;
      6'b000111 : _zz_shift_i_0_4 = shift_i_map_7;
      6'b001000 : _zz_shift_i_0_4 = shift_i_map_8;
      6'b001001 : _zz_shift_i_0_4 = shift_i_map_9;
      6'b001010 : _zz_shift_i_0_4 = shift_i_map_10;
      6'b001011 : _zz_shift_i_0_4 = shift_i_map_11;
      6'b001100 : _zz_shift_i_0_4 = shift_i_map_12;
      6'b001101 : _zz_shift_i_0_4 = shift_i_map_13;
      6'b001110 : _zz_shift_i_0_4 = shift_i_map_14;
      6'b001111 : _zz_shift_i_0_4 = shift_i_map_15;
      6'b010000 : _zz_shift_i_0_4 = shift_i_map_16;
      6'b010001 : _zz_shift_i_0_4 = shift_i_map_17;
      6'b010010 : _zz_shift_i_0_4 = shift_i_map_18;
      6'b010011 : _zz_shift_i_0_4 = shift_i_map_19;
      6'b010100 : _zz_shift_i_0_4 = shift_i_map_20;
      6'b010101 : _zz_shift_i_0_4 = shift_i_map_21;
      6'b010110 : _zz_shift_i_0_4 = shift_i_map_22;
      6'b010111 : _zz_shift_i_0_4 = shift_i_map_23;
      6'b011000 : _zz_shift_i_0_4 = shift_i_map_24;
      6'b011001 : _zz_shift_i_0_4 = shift_i_map_25;
      6'b011010 : _zz_shift_i_0_4 = shift_i_map_26;
      6'b011011 : _zz_shift_i_0_4 = shift_i_map_27;
      6'b011100 : _zz_shift_i_0_4 = shift_i_map_28;
      6'b011101 : _zz_shift_i_0_4 = shift_i_map_29;
      6'b011110 : _zz_shift_i_0_4 = shift_i_map_30;
      6'b011111 : _zz_shift_i_0_4 = shift_i_map_31;
      6'b100000 : _zz_shift_i_0_4 = shift_i_map_32;
      6'b100001 : _zz_shift_i_0_4 = shift_i_map_33;
      6'b100010 : _zz_shift_i_0_4 = shift_i_map_34;
      6'b100011 : _zz_shift_i_0_4 = shift_i_map_35;
      6'b100100 : _zz_shift_i_0_4 = shift_i_map_36;
      6'b100101 : _zz_shift_i_0_4 = shift_i_map_37;
      6'b100110 : _zz_shift_i_0_4 = shift_i_map_38;
      6'b100111 : _zz_shift_i_0_4 = shift_i_map_39;
      6'b101000 : _zz_shift_i_0_4 = shift_i_map_40;
      6'b101001 : _zz_shift_i_0_4 = shift_i_map_41;
      6'b101010 : _zz_shift_i_0_4 = shift_i_map_42;
      6'b101011 : _zz_shift_i_0_4 = shift_i_map_43;
      6'b101100 : _zz_shift_i_0_4 = shift_i_map_44;
      6'b101101 : _zz_shift_i_0_4 = shift_i_map_45;
      6'b101110 : _zz_shift_i_0_4 = shift_i_map_46;
      6'b101111 : _zz_shift_i_0_4 = shift_i_map_47;
      6'b110000 : _zz_shift_i_0_4 = shift_i_map_48;
      6'b110001 : _zz_shift_i_0_4 = shift_i_map_49;
      6'b110010 : _zz_shift_i_0_4 = shift_i_map_50;
      6'b110011 : _zz_shift_i_0_4 = shift_i_map_51;
      6'b110100 : _zz_shift_i_0_4 = shift_i_map_52;
      6'b110101 : _zz_shift_i_0_4 = shift_i_map_53;
      6'b110110 : _zz_shift_i_0_4 = shift_i_map_54;
      6'b110111 : _zz_shift_i_0_4 = shift_i_map_55;
      6'b111000 : _zz_shift_i_0_4 = shift_i_map_56;
      6'b111001 : _zz_shift_i_0_4 = shift_i_map_57;
      6'b111010 : _zz_shift_i_0_4 = shift_i_map_58;
      6'b111011 : _zz_shift_i_0_4 = shift_i_map_59;
      6'b111100 : _zz_shift_i_0_4 = shift_i_map_60;
      6'b111101 : _zz_shift_i_0_4 = shift_i_map_61;
      6'b111110 : _zz_shift_i_0_4 = shift_i_map_62;
      default : _zz_shift_i_0_4 = shift_i_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_0_5)
      6'b000000 : _zz_shift_q_0_4 = shift_q_map_0;
      6'b000001 : _zz_shift_q_0_4 = shift_q_map_1;
      6'b000010 : _zz_shift_q_0_4 = shift_q_map_2;
      6'b000011 : _zz_shift_q_0_4 = shift_q_map_3;
      6'b000100 : _zz_shift_q_0_4 = shift_q_map_4;
      6'b000101 : _zz_shift_q_0_4 = shift_q_map_5;
      6'b000110 : _zz_shift_q_0_4 = shift_q_map_6;
      6'b000111 : _zz_shift_q_0_4 = shift_q_map_7;
      6'b001000 : _zz_shift_q_0_4 = shift_q_map_8;
      6'b001001 : _zz_shift_q_0_4 = shift_q_map_9;
      6'b001010 : _zz_shift_q_0_4 = shift_q_map_10;
      6'b001011 : _zz_shift_q_0_4 = shift_q_map_11;
      6'b001100 : _zz_shift_q_0_4 = shift_q_map_12;
      6'b001101 : _zz_shift_q_0_4 = shift_q_map_13;
      6'b001110 : _zz_shift_q_0_4 = shift_q_map_14;
      6'b001111 : _zz_shift_q_0_4 = shift_q_map_15;
      6'b010000 : _zz_shift_q_0_4 = shift_q_map_16;
      6'b010001 : _zz_shift_q_0_4 = shift_q_map_17;
      6'b010010 : _zz_shift_q_0_4 = shift_q_map_18;
      6'b010011 : _zz_shift_q_0_4 = shift_q_map_19;
      6'b010100 : _zz_shift_q_0_4 = shift_q_map_20;
      6'b010101 : _zz_shift_q_0_4 = shift_q_map_21;
      6'b010110 : _zz_shift_q_0_4 = shift_q_map_22;
      6'b010111 : _zz_shift_q_0_4 = shift_q_map_23;
      6'b011000 : _zz_shift_q_0_4 = shift_q_map_24;
      6'b011001 : _zz_shift_q_0_4 = shift_q_map_25;
      6'b011010 : _zz_shift_q_0_4 = shift_q_map_26;
      6'b011011 : _zz_shift_q_0_4 = shift_q_map_27;
      6'b011100 : _zz_shift_q_0_4 = shift_q_map_28;
      6'b011101 : _zz_shift_q_0_4 = shift_q_map_29;
      6'b011110 : _zz_shift_q_0_4 = shift_q_map_30;
      6'b011111 : _zz_shift_q_0_4 = shift_q_map_31;
      6'b100000 : _zz_shift_q_0_4 = shift_q_map_32;
      6'b100001 : _zz_shift_q_0_4 = shift_q_map_33;
      6'b100010 : _zz_shift_q_0_4 = shift_q_map_34;
      6'b100011 : _zz_shift_q_0_4 = shift_q_map_35;
      6'b100100 : _zz_shift_q_0_4 = shift_q_map_36;
      6'b100101 : _zz_shift_q_0_4 = shift_q_map_37;
      6'b100110 : _zz_shift_q_0_4 = shift_q_map_38;
      6'b100111 : _zz_shift_q_0_4 = shift_q_map_39;
      6'b101000 : _zz_shift_q_0_4 = shift_q_map_40;
      6'b101001 : _zz_shift_q_0_4 = shift_q_map_41;
      6'b101010 : _zz_shift_q_0_4 = shift_q_map_42;
      6'b101011 : _zz_shift_q_0_4 = shift_q_map_43;
      6'b101100 : _zz_shift_q_0_4 = shift_q_map_44;
      6'b101101 : _zz_shift_q_0_4 = shift_q_map_45;
      6'b101110 : _zz_shift_q_0_4 = shift_q_map_46;
      6'b101111 : _zz_shift_q_0_4 = shift_q_map_47;
      6'b110000 : _zz_shift_q_0_4 = shift_q_map_48;
      6'b110001 : _zz_shift_q_0_4 = shift_q_map_49;
      6'b110010 : _zz_shift_q_0_4 = shift_q_map_50;
      6'b110011 : _zz_shift_q_0_4 = shift_q_map_51;
      6'b110100 : _zz_shift_q_0_4 = shift_q_map_52;
      6'b110101 : _zz_shift_q_0_4 = shift_q_map_53;
      6'b110110 : _zz_shift_q_0_4 = shift_q_map_54;
      6'b110111 : _zz_shift_q_0_4 = shift_q_map_55;
      6'b111000 : _zz_shift_q_0_4 = shift_q_map_56;
      6'b111001 : _zz_shift_q_0_4 = shift_q_map_57;
      6'b111010 : _zz_shift_q_0_4 = shift_q_map_58;
      6'b111011 : _zz_shift_q_0_4 = shift_q_map_59;
      6'b111100 : _zz_shift_q_0_4 = shift_q_map_60;
      6'b111101 : _zz_shift_q_0_4 = shift_q_map_61;
      6'b111110 : _zz_shift_q_0_4 = shift_q_map_62;
      default : _zz_shift_q_0_4 = shift_q_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_1_5)
      6'b000000 : _zz_shift_i_1_4 = shift_i_map_0;
      6'b000001 : _zz_shift_i_1_4 = shift_i_map_1;
      6'b000010 : _zz_shift_i_1_4 = shift_i_map_2;
      6'b000011 : _zz_shift_i_1_4 = shift_i_map_3;
      6'b000100 : _zz_shift_i_1_4 = shift_i_map_4;
      6'b000101 : _zz_shift_i_1_4 = shift_i_map_5;
      6'b000110 : _zz_shift_i_1_4 = shift_i_map_6;
      6'b000111 : _zz_shift_i_1_4 = shift_i_map_7;
      6'b001000 : _zz_shift_i_1_4 = shift_i_map_8;
      6'b001001 : _zz_shift_i_1_4 = shift_i_map_9;
      6'b001010 : _zz_shift_i_1_4 = shift_i_map_10;
      6'b001011 : _zz_shift_i_1_4 = shift_i_map_11;
      6'b001100 : _zz_shift_i_1_4 = shift_i_map_12;
      6'b001101 : _zz_shift_i_1_4 = shift_i_map_13;
      6'b001110 : _zz_shift_i_1_4 = shift_i_map_14;
      6'b001111 : _zz_shift_i_1_4 = shift_i_map_15;
      6'b010000 : _zz_shift_i_1_4 = shift_i_map_16;
      6'b010001 : _zz_shift_i_1_4 = shift_i_map_17;
      6'b010010 : _zz_shift_i_1_4 = shift_i_map_18;
      6'b010011 : _zz_shift_i_1_4 = shift_i_map_19;
      6'b010100 : _zz_shift_i_1_4 = shift_i_map_20;
      6'b010101 : _zz_shift_i_1_4 = shift_i_map_21;
      6'b010110 : _zz_shift_i_1_4 = shift_i_map_22;
      6'b010111 : _zz_shift_i_1_4 = shift_i_map_23;
      6'b011000 : _zz_shift_i_1_4 = shift_i_map_24;
      6'b011001 : _zz_shift_i_1_4 = shift_i_map_25;
      6'b011010 : _zz_shift_i_1_4 = shift_i_map_26;
      6'b011011 : _zz_shift_i_1_4 = shift_i_map_27;
      6'b011100 : _zz_shift_i_1_4 = shift_i_map_28;
      6'b011101 : _zz_shift_i_1_4 = shift_i_map_29;
      6'b011110 : _zz_shift_i_1_4 = shift_i_map_30;
      6'b011111 : _zz_shift_i_1_4 = shift_i_map_31;
      6'b100000 : _zz_shift_i_1_4 = shift_i_map_32;
      6'b100001 : _zz_shift_i_1_4 = shift_i_map_33;
      6'b100010 : _zz_shift_i_1_4 = shift_i_map_34;
      6'b100011 : _zz_shift_i_1_4 = shift_i_map_35;
      6'b100100 : _zz_shift_i_1_4 = shift_i_map_36;
      6'b100101 : _zz_shift_i_1_4 = shift_i_map_37;
      6'b100110 : _zz_shift_i_1_4 = shift_i_map_38;
      6'b100111 : _zz_shift_i_1_4 = shift_i_map_39;
      6'b101000 : _zz_shift_i_1_4 = shift_i_map_40;
      6'b101001 : _zz_shift_i_1_4 = shift_i_map_41;
      6'b101010 : _zz_shift_i_1_4 = shift_i_map_42;
      6'b101011 : _zz_shift_i_1_4 = shift_i_map_43;
      6'b101100 : _zz_shift_i_1_4 = shift_i_map_44;
      6'b101101 : _zz_shift_i_1_4 = shift_i_map_45;
      6'b101110 : _zz_shift_i_1_4 = shift_i_map_46;
      6'b101111 : _zz_shift_i_1_4 = shift_i_map_47;
      6'b110000 : _zz_shift_i_1_4 = shift_i_map_48;
      6'b110001 : _zz_shift_i_1_4 = shift_i_map_49;
      6'b110010 : _zz_shift_i_1_4 = shift_i_map_50;
      6'b110011 : _zz_shift_i_1_4 = shift_i_map_51;
      6'b110100 : _zz_shift_i_1_4 = shift_i_map_52;
      6'b110101 : _zz_shift_i_1_4 = shift_i_map_53;
      6'b110110 : _zz_shift_i_1_4 = shift_i_map_54;
      6'b110111 : _zz_shift_i_1_4 = shift_i_map_55;
      6'b111000 : _zz_shift_i_1_4 = shift_i_map_56;
      6'b111001 : _zz_shift_i_1_4 = shift_i_map_57;
      6'b111010 : _zz_shift_i_1_4 = shift_i_map_58;
      6'b111011 : _zz_shift_i_1_4 = shift_i_map_59;
      6'b111100 : _zz_shift_i_1_4 = shift_i_map_60;
      6'b111101 : _zz_shift_i_1_4 = shift_i_map_61;
      6'b111110 : _zz_shift_i_1_4 = shift_i_map_62;
      default : _zz_shift_i_1_4 = shift_i_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_1_5)
      6'b000000 : _zz_shift_q_1_4 = shift_q_map_0;
      6'b000001 : _zz_shift_q_1_4 = shift_q_map_1;
      6'b000010 : _zz_shift_q_1_4 = shift_q_map_2;
      6'b000011 : _zz_shift_q_1_4 = shift_q_map_3;
      6'b000100 : _zz_shift_q_1_4 = shift_q_map_4;
      6'b000101 : _zz_shift_q_1_4 = shift_q_map_5;
      6'b000110 : _zz_shift_q_1_4 = shift_q_map_6;
      6'b000111 : _zz_shift_q_1_4 = shift_q_map_7;
      6'b001000 : _zz_shift_q_1_4 = shift_q_map_8;
      6'b001001 : _zz_shift_q_1_4 = shift_q_map_9;
      6'b001010 : _zz_shift_q_1_4 = shift_q_map_10;
      6'b001011 : _zz_shift_q_1_4 = shift_q_map_11;
      6'b001100 : _zz_shift_q_1_4 = shift_q_map_12;
      6'b001101 : _zz_shift_q_1_4 = shift_q_map_13;
      6'b001110 : _zz_shift_q_1_4 = shift_q_map_14;
      6'b001111 : _zz_shift_q_1_4 = shift_q_map_15;
      6'b010000 : _zz_shift_q_1_4 = shift_q_map_16;
      6'b010001 : _zz_shift_q_1_4 = shift_q_map_17;
      6'b010010 : _zz_shift_q_1_4 = shift_q_map_18;
      6'b010011 : _zz_shift_q_1_4 = shift_q_map_19;
      6'b010100 : _zz_shift_q_1_4 = shift_q_map_20;
      6'b010101 : _zz_shift_q_1_4 = shift_q_map_21;
      6'b010110 : _zz_shift_q_1_4 = shift_q_map_22;
      6'b010111 : _zz_shift_q_1_4 = shift_q_map_23;
      6'b011000 : _zz_shift_q_1_4 = shift_q_map_24;
      6'b011001 : _zz_shift_q_1_4 = shift_q_map_25;
      6'b011010 : _zz_shift_q_1_4 = shift_q_map_26;
      6'b011011 : _zz_shift_q_1_4 = shift_q_map_27;
      6'b011100 : _zz_shift_q_1_4 = shift_q_map_28;
      6'b011101 : _zz_shift_q_1_4 = shift_q_map_29;
      6'b011110 : _zz_shift_q_1_4 = shift_q_map_30;
      6'b011111 : _zz_shift_q_1_4 = shift_q_map_31;
      6'b100000 : _zz_shift_q_1_4 = shift_q_map_32;
      6'b100001 : _zz_shift_q_1_4 = shift_q_map_33;
      6'b100010 : _zz_shift_q_1_4 = shift_q_map_34;
      6'b100011 : _zz_shift_q_1_4 = shift_q_map_35;
      6'b100100 : _zz_shift_q_1_4 = shift_q_map_36;
      6'b100101 : _zz_shift_q_1_4 = shift_q_map_37;
      6'b100110 : _zz_shift_q_1_4 = shift_q_map_38;
      6'b100111 : _zz_shift_q_1_4 = shift_q_map_39;
      6'b101000 : _zz_shift_q_1_4 = shift_q_map_40;
      6'b101001 : _zz_shift_q_1_4 = shift_q_map_41;
      6'b101010 : _zz_shift_q_1_4 = shift_q_map_42;
      6'b101011 : _zz_shift_q_1_4 = shift_q_map_43;
      6'b101100 : _zz_shift_q_1_4 = shift_q_map_44;
      6'b101101 : _zz_shift_q_1_4 = shift_q_map_45;
      6'b101110 : _zz_shift_q_1_4 = shift_q_map_46;
      6'b101111 : _zz_shift_q_1_4 = shift_q_map_47;
      6'b110000 : _zz_shift_q_1_4 = shift_q_map_48;
      6'b110001 : _zz_shift_q_1_4 = shift_q_map_49;
      6'b110010 : _zz_shift_q_1_4 = shift_q_map_50;
      6'b110011 : _zz_shift_q_1_4 = shift_q_map_51;
      6'b110100 : _zz_shift_q_1_4 = shift_q_map_52;
      6'b110101 : _zz_shift_q_1_4 = shift_q_map_53;
      6'b110110 : _zz_shift_q_1_4 = shift_q_map_54;
      6'b110111 : _zz_shift_q_1_4 = shift_q_map_55;
      6'b111000 : _zz_shift_q_1_4 = shift_q_map_56;
      6'b111001 : _zz_shift_q_1_4 = shift_q_map_57;
      6'b111010 : _zz_shift_q_1_4 = shift_q_map_58;
      6'b111011 : _zz_shift_q_1_4 = shift_q_map_59;
      6'b111100 : _zz_shift_q_1_4 = shift_q_map_60;
      6'b111101 : _zz_shift_q_1_4 = shift_q_map_61;
      6'b111110 : _zz_shift_q_1_4 = shift_q_map_62;
      default : _zz_shift_q_1_4 = shift_q_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_2_5)
      6'b000000 : _zz_shift_i_2_4 = shift_i_map_0;
      6'b000001 : _zz_shift_i_2_4 = shift_i_map_1;
      6'b000010 : _zz_shift_i_2_4 = shift_i_map_2;
      6'b000011 : _zz_shift_i_2_4 = shift_i_map_3;
      6'b000100 : _zz_shift_i_2_4 = shift_i_map_4;
      6'b000101 : _zz_shift_i_2_4 = shift_i_map_5;
      6'b000110 : _zz_shift_i_2_4 = shift_i_map_6;
      6'b000111 : _zz_shift_i_2_4 = shift_i_map_7;
      6'b001000 : _zz_shift_i_2_4 = shift_i_map_8;
      6'b001001 : _zz_shift_i_2_4 = shift_i_map_9;
      6'b001010 : _zz_shift_i_2_4 = shift_i_map_10;
      6'b001011 : _zz_shift_i_2_4 = shift_i_map_11;
      6'b001100 : _zz_shift_i_2_4 = shift_i_map_12;
      6'b001101 : _zz_shift_i_2_4 = shift_i_map_13;
      6'b001110 : _zz_shift_i_2_4 = shift_i_map_14;
      6'b001111 : _zz_shift_i_2_4 = shift_i_map_15;
      6'b010000 : _zz_shift_i_2_4 = shift_i_map_16;
      6'b010001 : _zz_shift_i_2_4 = shift_i_map_17;
      6'b010010 : _zz_shift_i_2_4 = shift_i_map_18;
      6'b010011 : _zz_shift_i_2_4 = shift_i_map_19;
      6'b010100 : _zz_shift_i_2_4 = shift_i_map_20;
      6'b010101 : _zz_shift_i_2_4 = shift_i_map_21;
      6'b010110 : _zz_shift_i_2_4 = shift_i_map_22;
      6'b010111 : _zz_shift_i_2_4 = shift_i_map_23;
      6'b011000 : _zz_shift_i_2_4 = shift_i_map_24;
      6'b011001 : _zz_shift_i_2_4 = shift_i_map_25;
      6'b011010 : _zz_shift_i_2_4 = shift_i_map_26;
      6'b011011 : _zz_shift_i_2_4 = shift_i_map_27;
      6'b011100 : _zz_shift_i_2_4 = shift_i_map_28;
      6'b011101 : _zz_shift_i_2_4 = shift_i_map_29;
      6'b011110 : _zz_shift_i_2_4 = shift_i_map_30;
      6'b011111 : _zz_shift_i_2_4 = shift_i_map_31;
      6'b100000 : _zz_shift_i_2_4 = shift_i_map_32;
      6'b100001 : _zz_shift_i_2_4 = shift_i_map_33;
      6'b100010 : _zz_shift_i_2_4 = shift_i_map_34;
      6'b100011 : _zz_shift_i_2_4 = shift_i_map_35;
      6'b100100 : _zz_shift_i_2_4 = shift_i_map_36;
      6'b100101 : _zz_shift_i_2_4 = shift_i_map_37;
      6'b100110 : _zz_shift_i_2_4 = shift_i_map_38;
      6'b100111 : _zz_shift_i_2_4 = shift_i_map_39;
      6'b101000 : _zz_shift_i_2_4 = shift_i_map_40;
      6'b101001 : _zz_shift_i_2_4 = shift_i_map_41;
      6'b101010 : _zz_shift_i_2_4 = shift_i_map_42;
      6'b101011 : _zz_shift_i_2_4 = shift_i_map_43;
      6'b101100 : _zz_shift_i_2_4 = shift_i_map_44;
      6'b101101 : _zz_shift_i_2_4 = shift_i_map_45;
      6'b101110 : _zz_shift_i_2_4 = shift_i_map_46;
      6'b101111 : _zz_shift_i_2_4 = shift_i_map_47;
      6'b110000 : _zz_shift_i_2_4 = shift_i_map_48;
      6'b110001 : _zz_shift_i_2_4 = shift_i_map_49;
      6'b110010 : _zz_shift_i_2_4 = shift_i_map_50;
      6'b110011 : _zz_shift_i_2_4 = shift_i_map_51;
      6'b110100 : _zz_shift_i_2_4 = shift_i_map_52;
      6'b110101 : _zz_shift_i_2_4 = shift_i_map_53;
      6'b110110 : _zz_shift_i_2_4 = shift_i_map_54;
      6'b110111 : _zz_shift_i_2_4 = shift_i_map_55;
      6'b111000 : _zz_shift_i_2_4 = shift_i_map_56;
      6'b111001 : _zz_shift_i_2_4 = shift_i_map_57;
      6'b111010 : _zz_shift_i_2_4 = shift_i_map_58;
      6'b111011 : _zz_shift_i_2_4 = shift_i_map_59;
      6'b111100 : _zz_shift_i_2_4 = shift_i_map_60;
      6'b111101 : _zz_shift_i_2_4 = shift_i_map_61;
      6'b111110 : _zz_shift_i_2_4 = shift_i_map_62;
      default : _zz_shift_i_2_4 = shift_i_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_2_5)
      6'b000000 : _zz_shift_q_2_4 = shift_q_map_0;
      6'b000001 : _zz_shift_q_2_4 = shift_q_map_1;
      6'b000010 : _zz_shift_q_2_4 = shift_q_map_2;
      6'b000011 : _zz_shift_q_2_4 = shift_q_map_3;
      6'b000100 : _zz_shift_q_2_4 = shift_q_map_4;
      6'b000101 : _zz_shift_q_2_4 = shift_q_map_5;
      6'b000110 : _zz_shift_q_2_4 = shift_q_map_6;
      6'b000111 : _zz_shift_q_2_4 = shift_q_map_7;
      6'b001000 : _zz_shift_q_2_4 = shift_q_map_8;
      6'b001001 : _zz_shift_q_2_4 = shift_q_map_9;
      6'b001010 : _zz_shift_q_2_4 = shift_q_map_10;
      6'b001011 : _zz_shift_q_2_4 = shift_q_map_11;
      6'b001100 : _zz_shift_q_2_4 = shift_q_map_12;
      6'b001101 : _zz_shift_q_2_4 = shift_q_map_13;
      6'b001110 : _zz_shift_q_2_4 = shift_q_map_14;
      6'b001111 : _zz_shift_q_2_4 = shift_q_map_15;
      6'b010000 : _zz_shift_q_2_4 = shift_q_map_16;
      6'b010001 : _zz_shift_q_2_4 = shift_q_map_17;
      6'b010010 : _zz_shift_q_2_4 = shift_q_map_18;
      6'b010011 : _zz_shift_q_2_4 = shift_q_map_19;
      6'b010100 : _zz_shift_q_2_4 = shift_q_map_20;
      6'b010101 : _zz_shift_q_2_4 = shift_q_map_21;
      6'b010110 : _zz_shift_q_2_4 = shift_q_map_22;
      6'b010111 : _zz_shift_q_2_4 = shift_q_map_23;
      6'b011000 : _zz_shift_q_2_4 = shift_q_map_24;
      6'b011001 : _zz_shift_q_2_4 = shift_q_map_25;
      6'b011010 : _zz_shift_q_2_4 = shift_q_map_26;
      6'b011011 : _zz_shift_q_2_4 = shift_q_map_27;
      6'b011100 : _zz_shift_q_2_4 = shift_q_map_28;
      6'b011101 : _zz_shift_q_2_4 = shift_q_map_29;
      6'b011110 : _zz_shift_q_2_4 = shift_q_map_30;
      6'b011111 : _zz_shift_q_2_4 = shift_q_map_31;
      6'b100000 : _zz_shift_q_2_4 = shift_q_map_32;
      6'b100001 : _zz_shift_q_2_4 = shift_q_map_33;
      6'b100010 : _zz_shift_q_2_4 = shift_q_map_34;
      6'b100011 : _zz_shift_q_2_4 = shift_q_map_35;
      6'b100100 : _zz_shift_q_2_4 = shift_q_map_36;
      6'b100101 : _zz_shift_q_2_4 = shift_q_map_37;
      6'b100110 : _zz_shift_q_2_4 = shift_q_map_38;
      6'b100111 : _zz_shift_q_2_4 = shift_q_map_39;
      6'b101000 : _zz_shift_q_2_4 = shift_q_map_40;
      6'b101001 : _zz_shift_q_2_4 = shift_q_map_41;
      6'b101010 : _zz_shift_q_2_4 = shift_q_map_42;
      6'b101011 : _zz_shift_q_2_4 = shift_q_map_43;
      6'b101100 : _zz_shift_q_2_4 = shift_q_map_44;
      6'b101101 : _zz_shift_q_2_4 = shift_q_map_45;
      6'b101110 : _zz_shift_q_2_4 = shift_q_map_46;
      6'b101111 : _zz_shift_q_2_4 = shift_q_map_47;
      6'b110000 : _zz_shift_q_2_4 = shift_q_map_48;
      6'b110001 : _zz_shift_q_2_4 = shift_q_map_49;
      6'b110010 : _zz_shift_q_2_4 = shift_q_map_50;
      6'b110011 : _zz_shift_q_2_4 = shift_q_map_51;
      6'b110100 : _zz_shift_q_2_4 = shift_q_map_52;
      6'b110101 : _zz_shift_q_2_4 = shift_q_map_53;
      6'b110110 : _zz_shift_q_2_4 = shift_q_map_54;
      6'b110111 : _zz_shift_q_2_4 = shift_q_map_55;
      6'b111000 : _zz_shift_q_2_4 = shift_q_map_56;
      6'b111001 : _zz_shift_q_2_4 = shift_q_map_57;
      6'b111010 : _zz_shift_q_2_4 = shift_q_map_58;
      6'b111011 : _zz_shift_q_2_4 = shift_q_map_59;
      6'b111100 : _zz_shift_q_2_4 = shift_q_map_60;
      6'b111101 : _zz_shift_q_2_4 = shift_q_map_61;
      6'b111110 : _zz_shift_q_2_4 = shift_q_map_62;
      default : _zz_shift_q_2_4 = shift_q_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_3_5)
      6'b000000 : _zz_shift_i_3_4 = shift_i_map_0;
      6'b000001 : _zz_shift_i_3_4 = shift_i_map_1;
      6'b000010 : _zz_shift_i_3_4 = shift_i_map_2;
      6'b000011 : _zz_shift_i_3_4 = shift_i_map_3;
      6'b000100 : _zz_shift_i_3_4 = shift_i_map_4;
      6'b000101 : _zz_shift_i_3_4 = shift_i_map_5;
      6'b000110 : _zz_shift_i_3_4 = shift_i_map_6;
      6'b000111 : _zz_shift_i_3_4 = shift_i_map_7;
      6'b001000 : _zz_shift_i_3_4 = shift_i_map_8;
      6'b001001 : _zz_shift_i_3_4 = shift_i_map_9;
      6'b001010 : _zz_shift_i_3_4 = shift_i_map_10;
      6'b001011 : _zz_shift_i_3_4 = shift_i_map_11;
      6'b001100 : _zz_shift_i_3_4 = shift_i_map_12;
      6'b001101 : _zz_shift_i_3_4 = shift_i_map_13;
      6'b001110 : _zz_shift_i_3_4 = shift_i_map_14;
      6'b001111 : _zz_shift_i_3_4 = shift_i_map_15;
      6'b010000 : _zz_shift_i_3_4 = shift_i_map_16;
      6'b010001 : _zz_shift_i_3_4 = shift_i_map_17;
      6'b010010 : _zz_shift_i_3_4 = shift_i_map_18;
      6'b010011 : _zz_shift_i_3_4 = shift_i_map_19;
      6'b010100 : _zz_shift_i_3_4 = shift_i_map_20;
      6'b010101 : _zz_shift_i_3_4 = shift_i_map_21;
      6'b010110 : _zz_shift_i_3_4 = shift_i_map_22;
      6'b010111 : _zz_shift_i_3_4 = shift_i_map_23;
      6'b011000 : _zz_shift_i_3_4 = shift_i_map_24;
      6'b011001 : _zz_shift_i_3_4 = shift_i_map_25;
      6'b011010 : _zz_shift_i_3_4 = shift_i_map_26;
      6'b011011 : _zz_shift_i_3_4 = shift_i_map_27;
      6'b011100 : _zz_shift_i_3_4 = shift_i_map_28;
      6'b011101 : _zz_shift_i_3_4 = shift_i_map_29;
      6'b011110 : _zz_shift_i_3_4 = shift_i_map_30;
      6'b011111 : _zz_shift_i_3_4 = shift_i_map_31;
      6'b100000 : _zz_shift_i_3_4 = shift_i_map_32;
      6'b100001 : _zz_shift_i_3_4 = shift_i_map_33;
      6'b100010 : _zz_shift_i_3_4 = shift_i_map_34;
      6'b100011 : _zz_shift_i_3_4 = shift_i_map_35;
      6'b100100 : _zz_shift_i_3_4 = shift_i_map_36;
      6'b100101 : _zz_shift_i_3_4 = shift_i_map_37;
      6'b100110 : _zz_shift_i_3_4 = shift_i_map_38;
      6'b100111 : _zz_shift_i_3_4 = shift_i_map_39;
      6'b101000 : _zz_shift_i_3_4 = shift_i_map_40;
      6'b101001 : _zz_shift_i_3_4 = shift_i_map_41;
      6'b101010 : _zz_shift_i_3_4 = shift_i_map_42;
      6'b101011 : _zz_shift_i_3_4 = shift_i_map_43;
      6'b101100 : _zz_shift_i_3_4 = shift_i_map_44;
      6'b101101 : _zz_shift_i_3_4 = shift_i_map_45;
      6'b101110 : _zz_shift_i_3_4 = shift_i_map_46;
      6'b101111 : _zz_shift_i_3_4 = shift_i_map_47;
      6'b110000 : _zz_shift_i_3_4 = shift_i_map_48;
      6'b110001 : _zz_shift_i_3_4 = shift_i_map_49;
      6'b110010 : _zz_shift_i_3_4 = shift_i_map_50;
      6'b110011 : _zz_shift_i_3_4 = shift_i_map_51;
      6'b110100 : _zz_shift_i_3_4 = shift_i_map_52;
      6'b110101 : _zz_shift_i_3_4 = shift_i_map_53;
      6'b110110 : _zz_shift_i_3_4 = shift_i_map_54;
      6'b110111 : _zz_shift_i_3_4 = shift_i_map_55;
      6'b111000 : _zz_shift_i_3_4 = shift_i_map_56;
      6'b111001 : _zz_shift_i_3_4 = shift_i_map_57;
      6'b111010 : _zz_shift_i_3_4 = shift_i_map_58;
      6'b111011 : _zz_shift_i_3_4 = shift_i_map_59;
      6'b111100 : _zz_shift_i_3_4 = shift_i_map_60;
      6'b111101 : _zz_shift_i_3_4 = shift_i_map_61;
      6'b111110 : _zz_shift_i_3_4 = shift_i_map_62;
      default : _zz_shift_i_3_4 = shift_i_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_3_5)
      6'b000000 : _zz_shift_q_3_4 = shift_q_map_0;
      6'b000001 : _zz_shift_q_3_4 = shift_q_map_1;
      6'b000010 : _zz_shift_q_3_4 = shift_q_map_2;
      6'b000011 : _zz_shift_q_3_4 = shift_q_map_3;
      6'b000100 : _zz_shift_q_3_4 = shift_q_map_4;
      6'b000101 : _zz_shift_q_3_4 = shift_q_map_5;
      6'b000110 : _zz_shift_q_3_4 = shift_q_map_6;
      6'b000111 : _zz_shift_q_3_4 = shift_q_map_7;
      6'b001000 : _zz_shift_q_3_4 = shift_q_map_8;
      6'b001001 : _zz_shift_q_3_4 = shift_q_map_9;
      6'b001010 : _zz_shift_q_3_4 = shift_q_map_10;
      6'b001011 : _zz_shift_q_3_4 = shift_q_map_11;
      6'b001100 : _zz_shift_q_3_4 = shift_q_map_12;
      6'b001101 : _zz_shift_q_3_4 = shift_q_map_13;
      6'b001110 : _zz_shift_q_3_4 = shift_q_map_14;
      6'b001111 : _zz_shift_q_3_4 = shift_q_map_15;
      6'b010000 : _zz_shift_q_3_4 = shift_q_map_16;
      6'b010001 : _zz_shift_q_3_4 = shift_q_map_17;
      6'b010010 : _zz_shift_q_3_4 = shift_q_map_18;
      6'b010011 : _zz_shift_q_3_4 = shift_q_map_19;
      6'b010100 : _zz_shift_q_3_4 = shift_q_map_20;
      6'b010101 : _zz_shift_q_3_4 = shift_q_map_21;
      6'b010110 : _zz_shift_q_3_4 = shift_q_map_22;
      6'b010111 : _zz_shift_q_3_4 = shift_q_map_23;
      6'b011000 : _zz_shift_q_3_4 = shift_q_map_24;
      6'b011001 : _zz_shift_q_3_4 = shift_q_map_25;
      6'b011010 : _zz_shift_q_3_4 = shift_q_map_26;
      6'b011011 : _zz_shift_q_3_4 = shift_q_map_27;
      6'b011100 : _zz_shift_q_3_4 = shift_q_map_28;
      6'b011101 : _zz_shift_q_3_4 = shift_q_map_29;
      6'b011110 : _zz_shift_q_3_4 = shift_q_map_30;
      6'b011111 : _zz_shift_q_3_4 = shift_q_map_31;
      6'b100000 : _zz_shift_q_3_4 = shift_q_map_32;
      6'b100001 : _zz_shift_q_3_4 = shift_q_map_33;
      6'b100010 : _zz_shift_q_3_4 = shift_q_map_34;
      6'b100011 : _zz_shift_q_3_4 = shift_q_map_35;
      6'b100100 : _zz_shift_q_3_4 = shift_q_map_36;
      6'b100101 : _zz_shift_q_3_4 = shift_q_map_37;
      6'b100110 : _zz_shift_q_3_4 = shift_q_map_38;
      6'b100111 : _zz_shift_q_3_4 = shift_q_map_39;
      6'b101000 : _zz_shift_q_3_4 = shift_q_map_40;
      6'b101001 : _zz_shift_q_3_4 = shift_q_map_41;
      6'b101010 : _zz_shift_q_3_4 = shift_q_map_42;
      6'b101011 : _zz_shift_q_3_4 = shift_q_map_43;
      6'b101100 : _zz_shift_q_3_4 = shift_q_map_44;
      6'b101101 : _zz_shift_q_3_4 = shift_q_map_45;
      6'b101110 : _zz_shift_q_3_4 = shift_q_map_46;
      6'b101111 : _zz_shift_q_3_4 = shift_q_map_47;
      6'b110000 : _zz_shift_q_3_4 = shift_q_map_48;
      6'b110001 : _zz_shift_q_3_4 = shift_q_map_49;
      6'b110010 : _zz_shift_q_3_4 = shift_q_map_50;
      6'b110011 : _zz_shift_q_3_4 = shift_q_map_51;
      6'b110100 : _zz_shift_q_3_4 = shift_q_map_52;
      6'b110101 : _zz_shift_q_3_4 = shift_q_map_53;
      6'b110110 : _zz_shift_q_3_4 = shift_q_map_54;
      6'b110111 : _zz_shift_q_3_4 = shift_q_map_55;
      6'b111000 : _zz_shift_q_3_4 = shift_q_map_56;
      6'b111001 : _zz_shift_q_3_4 = shift_q_map_57;
      6'b111010 : _zz_shift_q_3_4 = shift_q_map_58;
      6'b111011 : _zz_shift_q_3_4 = shift_q_map_59;
      6'b111100 : _zz_shift_q_3_4 = shift_q_map_60;
      6'b111101 : _zz_shift_q_3_4 = shift_q_map_61;
      6'b111110 : _zz_shift_q_3_4 = shift_q_map_62;
      default : _zz_shift_q_3_4 = shift_q_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_4_5)
      6'b000000 : _zz_shift_i_4_4 = shift_i_map_0;
      6'b000001 : _zz_shift_i_4_4 = shift_i_map_1;
      6'b000010 : _zz_shift_i_4_4 = shift_i_map_2;
      6'b000011 : _zz_shift_i_4_4 = shift_i_map_3;
      6'b000100 : _zz_shift_i_4_4 = shift_i_map_4;
      6'b000101 : _zz_shift_i_4_4 = shift_i_map_5;
      6'b000110 : _zz_shift_i_4_4 = shift_i_map_6;
      6'b000111 : _zz_shift_i_4_4 = shift_i_map_7;
      6'b001000 : _zz_shift_i_4_4 = shift_i_map_8;
      6'b001001 : _zz_shift_i_4_4 = shift_i_map_9;
      6'b001010 : _zz_shift_i_4_4 = shift_i_map_10;
      6'b001011 : _zz_shift_i_4_4 = shift_i_map_11;
      6'b001100 : _zz_shift_i_4_4 = shift_i_map_12;
      6'b001101 : _zz_shift_i_4_4 = shift_i_map_13;
      6'b001110 : _zz_shift_i_4_4 = shift_i_map_14;
      6'b001111 : _zz_shift_i_4_4 = shift_i_map_15;
      6'b010000 : _zz_shift_i_4_4 = shift_i_map_16;
      6'b010001 : _zz_shift_i_4_4 = shift_i_map_17;
      6'b010010 : _zz_shift_i_4_4 = shift_i_map_18;
      6'b010011 : _zz_shift_i_4_4 = shift_i_map_19;
      6'b010100 : _zz_shift_i_4_4 = shift_i_map_20;
      6'b010101 : _zz_shift_i_4_4 = shift_i_map_21;
      6'b010110 : _zz_shift_i_4_4 = shift_i_map_22;
      6'b010111 : _zz_shift_i_4_4 = shift_i_map_23;
      6'b011000 : _zz_shift_i_4_4 = shift_i_map_24;
      6'b011001 : _zz_shift_i_4_4 = shift_i_map_25;
      6'b011010 : _zz_shift_i_4_4 = shift_i_map_26;
      6'b011011 : _zz_shift_i_4_4 = shift_i_map_27;
      6'b011100 : _zz_shift_i_4_4 = shift_i_map_28;
      6'b011101 : _zz_shift_i_4_4 = shift_i_map_29;
      6'b011110 : _zz_shift_i_4_4 = shift_i_map_30;
      6'b011111 : _zz_shift_i_4_4 = shift_i_map_31;
      6'b100000 : _zz_shift_i_4_4 = shift_i_map_32;
      6'b100001 : _zz_shift_i_4_4 = shift_i_map_33;
      6'b100010 : _zz_shift_i_4_4 = shift_i_map_34;
      6'b100011 : _zz_shift_i_4_4 = shift_i_map_35;
      6'b100100 : _zz_shift_i_4_4 = shift_i_map_36;
      6'b100101 : _zz_shift_i_4_4 = shift_i_map_37;
      6'b100110 : _zz_shift_i_4_4 = shift_i_map_38;
      6'b100111 : _zz_shift_i_4_4 = shift_i_map_39;
      6'b101000 : _zz_shift_i_4_4 = shift_i_map_40;
      6'b101001 : _zz_shift_i_4_4 = shift_i_map_41;
      6'b101010 : _zz_shift_i_4_4 = shift_i_map_42;
      6'b101011 : _zz_shift_i_4_4 = shift_i_map_43;
      6'b101100 : _zz_shift_i_4_4 = shift_i_map_44;
      6'b101101 : _zz_shift_i_4_4 = shift_i_map_45;
      6'b101110 : _zz_shift_i_4_4 = shift_i_map_46;
      6'b101111 : _zz_shift_i_4_4 = shift_i_map_47;
      6'b110000 : _zz_shift_i_4_4 = shift_i_map_48;
      6'b110001 : _zz_shift_i_4_4 = shift_i_map_49;
      6'b110010 : _zz_shift_i_4_4 = shift_i_map_50;
      6'b110011 : _zz_shift_i_4_4 = shift_i_map_51;
      6'b110100 : _zz_shift_i_4_4 = shift_i_map_52;
      6'b110101 : _zz_shift_i_4_4 = shift_i_map_53;
      6'b110110 : _zz_shift_i_4_4 = shift_i_map_54;
      6'b110111 : _zz_shift_i_4_4 = shift_i_map_55;
      6'b111000 : _zz_shift_i_4_4 = shift_i_map_56;
      6'b111001 : _zz_shift_i_4_4 = shift_i_map_57;
      6'b111010 : _zz_shift_i_4_4 = shift_i_map_58;
      6'b111011 : _zz_shift_i_4_4 = shift_i_map_59;
      6'b111100 : _zz_shift_i_4_4 = shift_i_map_60;
      6'b111101 : _zz_shift_i_4_4 = shift_i_map_61;
      6'b111110 : _zz_shift_i_4_4 = shift_i_map_62;
      default : _zz_shift_i_4_4 = shift_i_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_4_5)
      6'b000000 : _zz_shift_q_4_4 = shift_q_map_0;
      6'b000001 : _zz_shift_q_4_4 = shift_q_map_1;
      6'b000010 : _zz_shift_q_4_4 = shift_q_map_2;
      6'b000011 : _zz_shift_q_4_4 = shift_q_map_3;
      6'b000100 : _zz_shift_q_4_4 = shift_q_map_4;
      6'b000101 : _zz_shift_q_4_4 = shift_q_map_5;
      6'b000110 : _zz_shift_q_4_4 = shift_q_map_6;
      6'b000111 : _zz_shift_q_4_4 = shift_q_map_7;
      6'b001000 : _zz_shift_q_4_4 = shift_q_map_8;
      6'b001001 : _zz_shift_q_4_4 = shift_q_map_9;
      6'b001010 : _zz_shift_q_4_4 = shift_q_map_10;
      6'b001011 : _zz_shift_q_4_4 = shift_q_map_11;
      6'b001100 : _zz_shift_q_4_4 = shift_q_map_12;
      6'b001101 : _zz_shift_q_4_4 = shift_q_map_13;
      6'b001110 : _zz_shift_q_4_4 = shift_q_map_14;
      6'b001111 : _zz_shift_q_4_4 = shift_q_map_15;
      6'b010000 : _zz_shift_q_4_4 = shift_q_map_16;
      6'b010001 : _zz_shift_q_4_4 = shift_q_map_17;
      6'b010010 : _zz_shift_q_4_4 = shift_q_map_18;
      6'b010011 : _zz_shift_q_4_4 = shift_q_map_19;
      6'b010100 : _zz_shift_q_4_4 = shift_q_map_20;
      6'b010101 : _zz_shift_q_4_4 = shift_q_map_21;
      6'b010110 : _zz_shift_q_4_4 = shift_q_map_22;
      6'b010111 : _zz_shift_q_4_4 = shift_q_map_23;
      6'b011000 : _zz_shift_q_4_4 = shift_q_map_24;
      6'b011001 : _zz_shift_q_4_4 = shift_q_map_25;
      6'b011010 : _zz_shift_q_4_4 = shift_q_map_26;
      6'b011011 : _zz_shift_q_4_4 = shift_q_map_27;
      6'b011100 : _zz_shift_q_4_4 = shift_q_map_28;
      6'b011101 : _zz_shift_q_4_4 = shift_q_map_29;
      6'b011110 : _zz_shift_q_4_4 = shift_q_map_30;
      6'b011111 : _zz_shift_q_4_4 = shift_q_map_31;
      6'b100000 : _zz_shift_q_4_4 = shift_q_map_32;
      6'b100001 : _zz_shift_q_4_4 = shift_q_map_33;
      6'b100010 : _zz_shift_q_4_4 = shift_q_map_34;
      6'b100011 : _zz_shift_q_4_4 = shift_q_map_35;
      6'b100100 : _zz_shift_q_4_4 = shift_q_map_36;
      6'b100101 : _zz_shift_q_4_4 = shift_q_map_37;
      6'b100110 : _zz_shift_q_4_4 = shift_q_map_38;
      6'b100111 : _zz_shift_q_4_4 = shift_q_map_39;
      6'b101000 : _zz_shift_q_4_4 = shift_q_map_40;
      6'b101001 : _zz_shift_q_4_4 = shift_q_map_41;
      6'b101010 : _zz_shift_q_4_4 = shift_q_map_42;
      6'b101011 : _zz_shift_q_4_4 = shift_q_map_43;
      6'b101100 : _zz_shift_q_4_4 = shift_q_map_44;
      6'b101101 : _zz_shift_q_4_4 = shift_q_map_45;
      6'b101110 : _zz_shift_q_4_4 = shift_q_map_46;
      6'b101111 : _zz_shift_q_4_4 = shift_q_map_47;
      6'b110000 : _zz_shift_q_4_4 = shift_q_map_48;
      6'b110001 : _zz_shift_q_4_4 = shift_q_map_49;
      6'b110010 : _zz_shift_q_4_4 = shift_q_map_50;
      6'b110011 : _zz_shift_q_4_4 = shift_q_map_51;
      6'b110100 : _zz_shift_q_4_4 = shift_q_map_52;
      6'b110101 : _zz_shift_q_4_4 = shift_q_map_53;
      6'b110110 : _zz_shift_q_4_4 = shift_q_map_54;
      6'b110111 : _zz_shift_q_4_4 = shift_q_map_55;
      6'b111000 : _zz_shift_q_4_4 = shift_q_map_56;
      6'b111001 : _zz_shift_q_4_4 = shift_q_map_57;
      6'b111010 : _zz_shift_q_4_4 = shift_q_map_58;
      6'b111011 : _zz_shift_q_4_4 = shift_q_map_59;
      6'b111100 : _zz_shift_q_4_4 = shift_q_map_60;
      6'b111101 : _zz_shift_q_4_4 = shift_q_map_61;
      6'b111110 : _zz_shift_q_4_4 = shift_q_map_62;
      default : _zz_shift_q_4_4 = shift_q_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_5_5)
      6'b000000 : _zz_shift_i_5_4 = shift_i_map_0;
      6'b000001 : _zz_shift_i_5_4 = shift_i_map_1;
      6'b000010 : _zz_shift_i_5_4 = shift_i_map_2;
      6'b000011 : _zz_shift_i_5_4 = shift_i_map_3;
      6'b000100 : _zz_shift_i_5_4 = shift_i_map_4;
      6'b000101 : _zz_shift_i_5_4 = shift_i_map_5;
      6'b000110 : _zz_shift_i_5_4 = shift_i_map_6;
      6'b000111 : _zz_shift_i_5_4 = shift_i_map_7;
      6'b001000 : _zz_shift_i_5_4 = shift_i_map_8;
      6'b001001 : _zz_shift_i_5_4 = shift_i_map_9;
      6'b001010 : _zz_shift_i_5_4 = shift_i_map_10;
      6'b001011 : _zz_shift_i_5_4 = shift_i_map_11;
      6'b001100 : _zz_shift_i_5_4 = shift_i_map_12;
      6'b001101 : _zz_shift_i_5_4 = shift_i_map_13;
      6'b001110 : _zz_shift_i_5_4 = shift_i_map_14;
      6'b001111 : _zz_shift_i_5_4 = shift_i_map_15;
      6'b010000 : _zz_shift_i_5_4 = shift_i_map_16;
      6'b010001 : _zz_shift_i_5_4 = shift_i_map_17;
      6'b010010 : _zz_shift_i_5_4 = shift_i_map_18;
      6'b010011 : _zz_shift_i_5_4 = shift_i_map_19;
      6'b010100 : _zz_shift_i_5_4 = shift_i_map_20;
      6'b010101 : _zz_shift_i_5_4 = shift_i_map_21;
      6'b010110 : _zz_shift_i_5_4 = shift_i_map_22;
      6'b010111 : _zz_shift_i_5_4 = shift_i_map_23;
      6'b011000 : _zz_shift_i_5_4 = shift_i_map_24;
      6'b011001 : _zz_shift_i_5_4 = shift_i_map_25;
      6'b011010 : _zz_shift_i_5_4 = shift_i_map_26;
      6'b011011 : _zz_shift_i_5_4 = shift_i_map_27;
      6'b011100 : _zz_shift_i_5_4 = shift_i_map_28;
      6'b011101 : _zz_shift_i_5_4 = shift_i_map_29;
      6'b011110 : _zz_shift_i_5_4 = shift_i_map_30;
      6'b011111 : _zz_shift_i_5_4 = shift_i_map_31;
      6'b100000 : _zz_shift_i_5_4 = shift_i_map_32;
      6'b100001 : _zz_shift_i_5_4 = shift_i_map_33;
      6'b100010 : _zz_shift_i_5_4 = shift_i_map_34;
      6'b100011 : _zz_shift_i_5_4 = shift_i_map_35;
      6'b100100 : _zz_shift_i_5_4 = shift_i_map_36;
      6'b100101 : _zz_shift_i_5_4 = shift_i_map_37;
      6'b100110 : _zz_shift_i_5_4 = shift_i_map_38;
      6'b100111 : _zz_shift_i_5_4 = shift_i_map_39;
      6'b101000 : _zz_shift_i_5_4 = shift_i_map_40;
      6'b101001 : _zz_shift_i_5_4 = shift_i_map_41;
      6'b101010 : _zz_shift_i_5_4 = shift_i_map_42;
      6'b101011 : _zz_shift_i_5_4 = shift_i_map_43;
      6'b101100 : _zz_shift_i_5_4 = shift_i_map_44;
      6'b101101 : _zz_shift_i_5_4 = shift_i_map_45;
      6'b101110 : _zz_shift_i_5_4 = shift_i_map_46;
      6'b101111 : _zz_shift_i_5_4 = shift_i_map_47;
      6'b110000 : _zz_shift_i_5_4 = shift_i_map_48;
      6'b110001 : _zz_shift_i_5_4 = shift_i_map_49;
      6'b110010 : _zz_shift_i_5_4 = shift_i_map_50;
      6'b110011 : _zz_shift_i_5_4 = shift_i_map_51;
      6'b110100 : _zz_shift_i_5_4 = shift_i_map_52;
      6'b110101 : _zz_shift_i_5_4 = shift_i_map_53;
      6'b110110 : _zz_shift_i_5_4 = shift_i_map_54;
      6'b110111 : _zz_shift_i_5_4 = shift_i_map_55;
      6'b111000 : _zz_shift_i_5_4 = shift_i_map_56;
      6'b111001 : _zz_shift_i_5_4 = shift_i_map_57;
      6'b111010 : _zz_shift_i_5_4 = shift_i_map_58;
      6'b111011 : _zz_shift_i_5_4 = shift_i_map_59;
      6'b111100 : _zz_shift_i_5_4 = shift_i_map_60;
      6'b111101 : _zz_shift_i_5_4 = shift_i_map_61;
      6'b111110 : _zz_shift_i_5_4 = shift_i_map_62;
      default : _zz_shift_i_5_4 = shift_i_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_5_5)
      6'b000000 : _zz_shift_q_5_4 = shift_q_map_0;
      6'b000001 : _zz_shift_q_5_4 = shift_q_map_1;
      6'b000010 : _zz_shift_q_5_4 = shift_q_map_2;
      6'b000011 : _zz_shift_q_5_4 = shift_q_map_3;
      6'b000100 : _zz_shift_q_5_4 = shift_q_map_4;
      6'b000101 : _zz_shift_q_5_4 = shift_q_map_5;
      6'b000110 : _zz_shift_q_5_4 = shift_q_map_6;
      6'b000111 : _zz_shift_q_5_4 = shift_q_map_7;
      6'b001000 : _zz_shift_q_5_4 = shift_q_map_8;
      6'b001001 : _zz_shift_q_5_4 = shift_q_map_9;
      6'b001010 : _zz_shift_q_5_4 = shift_q_map_10;
      6'b001011 : _zz_shift_q_5_4 = shift_q_map_11;
      6'b001100 : _zz_shift_q_5_4 = shift_q_map_12;
      6'b001101 : _zz_shift_q_5_4 = shift_q_map_13;
      6'b001110 : _zz_shift_q_5_4 = shift_q_map_14;
      6'b001111 : _zz_shift_q_5_4 = shift_q_map_15;
      6'b010000 : _zz_shift_q_5_4 = shift_q_map_16;
      6'b010001 : _zz_shift_q_5_4 = shift_q_map_17;
      6'b010010 : _zz_shift_q_5_4 = shift_q_map_18;
      6'b010011 : _zz_shift_q_5_4 = shift_q_map_19;
      6'b010100 : _zz_shift_q_5_4 = shift_q_map_20;
      6'b010101 : _zz_shift_q_5_4 = shift_q_map_21;
      6'b010110 : _zz_shift_q_5_4 = shift_q_map_22;
      6'b010111 : _zz_shift_q_5_4 = shift_q_map_23;
      6'b011000 : _zz_shift_q_5_4 = shift_q_map_24;
      6'b011001 : _zz_shift_q_5_4 = shift_q_map_25;
      6'b011010 : _zz_shift_q_5_4 = shift_q_map_26;
      6'b011011 : _zz_shift_q_5_4 = shift_q_map_27;
      6'b011100 : _zz_shift_q_5_4 = shift_q_map_28;
      6'b011101 : _zz_shift_q_5_4 = shift_q_map_29;
      6'b011110 : _zz_shift_q_5_4 = shift_q_map_30;
      6'b011111 : _zz_shift_q_5_4 = shift_q_map_31;
      6'b100000 : _zz_shift_q_5_4 = shift_q_map_32;
      6'b100001 : _zz_shift_q_5_4 = shift_q_map_33;
      6'b100010 : _zz_shift_q_5_4 = shift_q_map_34;
      6'b100011 : _zz_shift_q_5_4 = shift_q_map_35;
      6'b100100 : _zz_shift_q_5_4 = shift_q_map_36;
      6'b100101 : _zz_shift_q_5_4 = shift_q_map_37;
      6'b100110 : _zz_shift_q_5_4 = shift_q_map_38;
      6'b100111 : _zz_shift_q_5_4 = shift_q_map_39;
      6'b101000 : _zz_shift_q_5_4 = shift_q_map_40;
      6'b101001 : _zz_shift_q_5_4 = shift_q_map_41;
      6'b101010 : _zz_shift_q_5_4 = shift_q_map_42;
      6'b101011 : _zz_shift_q_5_4 = shift_q_map_43;
      6'b101100 : _zz_shift_q_5_4 = shift_q_map_44;
      6'b101101 : _zz_shift_q_5_4 = shift_q_map_45;
      6'b101110 : _zz_shift_q_5_4 = shift_q_map_46;
      6'b101111 : _zz_shift_q_5_4 = shift_q_map_47;
      6'b110000 : _zz_shift_q_5_4 = shift_q_map_48;
      6'b110001 : _zz_shift_q_5_4 = shift_q_map_49;
      6'b110010 : _zz_shift_q_5_4 = shift_q_map_50;
      6'b110011 : _zz_shift_q_5_4 = shift_q_map_51;
      6'b110100 : _zz_shift_q_5_4 = shift_q_map_52;
      6'b110101 : _zz_shift_q_5_4 = shift_q_map_53;
      6'b110110 : _zz_shift_q_5_4 = shift_q_map_54;
      6'b110111 : _zz_shift_q_5_4 = shift_q_map_55;
      6'b111000 : _zz_shift_q_5_4 = shift_q_map_56;
      6'b111001 : _zz_shift_q_5_4 = shift_q_map_57;
      6'b111010 : _zz_shift_q_5_4 = shift_q_map_58;
      6'b111011 : _zz_shift_q_5_4 = shift_q_map_59;
      6'b111100 : _zz_shift_q_5_4 = shift_q_map_60;
      6'b111101 : _zz_shift_q_5_4 = shift_q_map_61;
      6'b111110 : _zz_shift_q_5_4 = shift_q_map_62;
      default : _zz_shift_q_5_4 = shift_q_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_6_5)
      6'b000000 : _zz_shift_i_6_4 = shift_i_map_0;
      6'b000001 : _zz_shift_i_6_4 = shift_i_map_1;
      6'b000010 : _zz_shift_i_6_4 = shift_i_map_2;
      6'b000011 : _zz_shift_i_6_4 = shift_i_map_3;
      6'b000100 : _zz_shift_i_6_4 = shift_i_map_4;
      6'b000101 : _zz_shift_i_6_4 = shift_i_map_5;
      6'b000110 : _zz_shift_i_6_4 = shift_i_map_6;
      6'b000111 : _zz_shift_i_6_4 = shift_i_map_7;
      6'b001000 : _zz_shift_i_6_4 = shift_i_map_8;
      6'b001001 : _zz_shift_i_6_4 = shift_i_map_9;
      6'b001010 : _zz_shift_i_6_4 = shift_i_map_10;
      6'b001011 : _zz_shift_i_6_4 = shift_i_map_11;
      6'b001100 : _zz_shift_i_6_4 = shift_i_map_12;
      6'b001101 : _zz_shift_i_6_4 = shift_i_map_13;
      6'b001110 : _zz_shift_i_6_4 = shift_i_map_14;
      6'b001111 : _zz_shift_i_6_4 = shift_i_map_15;
      6'b010000 : _zz_shift_i_6_4 = shift_i_map_16;
      6'b010001 : _zz_shift_i_6_4 = shift_i_map_17;
      6'b010010 : _zz_shift_i_6_4 = shift_i_map_18;
      6'b010011 : _zz_shift_i_6_4 = shift_i_map_19;
      6'b010100 : _zz_shift_i_6_4 = shift_i_map_20;
      6'b010101 : _zz_shift_i_6_4 = shift_i_map_21;
      6'b010110 : _zz_shift_i_6_4 = shift_i_map_22;
      6'b010111 : _zz_shift_i_6_4 = shift_i_map_23;
      6'b011000 : _zz_shift_i_6_4 = shift_i_map_24;
      6'b011001 : _zz_shift_i_6_4 = shift_i_map_25;
      6'b011010 : _zz_shift_i_6_4 = shift_i_map_26;
      6'b011011 : _zz_shift_i_6_4 = shift_i_map_27;
      6'b011100 : _zz_shift_i_6_4 = shift_i_map_28;
      6'b011101 : _zz_shift_i_6_4 = shift_i_map_29;
      6'b011110 : _zz_shift_i_6_4 = shift_i_map_30;
      6'b011111 : _zz_shift_i_6_4 = shift_i_map_31;
      6'b100000 : _zz_shift_i_6_4 = shift_i_map_32;
      6'b100001 : _zz_shift_i_6_4 = shift_i_map_33;
      6'b100010 : _zz_shift_i_6_4 = shift_i_map_34;
      6'b100011 : _zz_shift_i_6_4 = shift_i_map_35;
      6'b100100 : _zz_shift_i_6_4 = shift_i_map_36;
      6'b100101 : _zz_shift_i_6_4 = shift_i_map_37;
      6'b100110 : _zz_shift_i_6_4 = shift_i_map_38;
      6'b100111 : _zz_shift_i_6_4 = shift_i_map_39;
      6'b101000 : _zz_shift_i_6_4 = shift_i_map_40;
      6'b101001 : _zz_shift_i_6_4 = shift_i_map_41;
      6'b101010 : _zz_shift_i_6_4 = shift_i_map_42;
      6'b101011 : _zz_shift_i_6_4 = shift_i_map_43;
      6'b101100 : _zz_shift_i_6_4 = shift_i_map_44;
      6'b101101 : _zz_shift_i_6_4 = shift_i_map_45;
      6'b101110 : _zz_shift_i_6_4 = shift_i_map_46;
      6'b101111 : _zz_shift_i_6_4 = shift_i_map_47;
      6'b110000 : _zz_shift_i_6_4 = shift_i_map_48;
      6'b110001 : _zz_shift_i_6_4 = shift_i_map_49;
      6'b110010 : _zz_shift_i_6_4 = shift_i_map_50;
      6'b110011 : _zz_shift_i_6_4 = shift_i_map_51;
      6'b110100 : _zz_shift_i_6_4 = shift_i_map_52;
      6'b110101 : _zz_shift_i_6_4 = shift_i_map_53;
      6'b110110 : _zz_shift_i_6_4 = shift_i_map_54;
      6'b110111 : _zz_shift_i_6_4 = shift_i_map_55;
      6'b111000 : _zz_shift_i_6_4 = shift_i_map_56;
      6'b111001 : _zz_shift_i_6_4 = shift_i_map_57;
      6'b111010 : _zz_shift_i_6_4 = shift_i_map_58;
      6'b111011 : _zz_shift_i_6_4 = shift_i_map_59;
      6'b111100 : _zz_shift_i_6_4 = shift_i_map_60;
      6'b111101 : _zz_shift_i_6_4 = shift_i_map_61;
      6'b111110 : _zz_shift_i_6_4 = shift_i_map_62;
      default : _zz_shift_i_6_4 = shift_i_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_6_5)
      6'b000000 : _zz_shift_q_6_4 = shift_q_map_0;
      6'b000001 : _zz_shift_q_6_4 = shift_q_map_1;
      6'b000010 : _zz_shift_q_6_4 = shift_q_map_2;
      6'b000011 : _zz_shift_q_6_4 = shift_q_map_3;
      6'b000100 : _zz_shift_q_6_4 = shift_q_map_4;
      6'b000101 : _zz_shift_q_6_4 = shift_q_map_5;
      6'b000110 : _zz_shift_q_6_4 = shift_q_map_6;
      6'b000111 : _zz_shift_q_6_4 = shift_q_map_7;
      6'b001000 : _zz_shift_q_6_4 = shift_q_map_8;
      6'b001001 : _zz_shift_q_6_4 = shift_q_map_9;
      6'b001010 : _zz_shift_q_6_4 = shift_q_map_10;
      6'b001011 : _zz_shift_q_6_4 = shift_q_map_11;
      6'b001100 : _zz_shift_q_6_4 = shift_q_map_12;
      6'b001101 : _zz_shift_q_6_4 = shift_q_map_13;
      6'b001110 : _zz_shift_q_6_4 = shift_q_map_14;
      6'b001111 : _zz_shift_q_6_4 = shift_q_map_15;
      6'b010000 : _zz_shift_q_6_4 = shift_q_map_16;
      6'b010001 : _zz_shift_q_6_4 = shift_q_map_17;
      6'b010010 : _zz_shift_q_6_4 = shift_q_map_18;
      6'b010011 : _zz_shift_q_6_4 = shift_q_map_19;
      6'b010100 : _zz_shift_q_6_4 = shift_q_map_20;
      6'b010101 : _zz_shift_q_6_4 = shift_q_map_21;
      6'b010110 : _zz_shift_q_6_4 = shift_q_map_22;
      6'b010111 : _zz_shift_q_6_4 = shift_q_map_23;
      6'b011000 : _zz_shift_q_6_4 = shift_q_map_24;
      6'b011001 : _zz_shift_q_6_4 = shift_q_map_25;
      6'b011010 : _zz_shift_q_6_4 = shift_q_map_26;
      6'b011011 : _zz_shift_q_6_4 = shift_q_map_27;
      6'b011100 : _zz_shift_q_6_4 = shift_q_map_28;
      6'b011101 : _zz_shift_q_6_4 = shift_q_map_29;
      6'b011110 : _zz_shift_q_6_4 = shift_q_map_30;
      6'b011111 : _zz_shift_q_6_4 = shift_q_map_31;
      6'b100000 : _zz_shift_q_6_4 = shift_q_map_32;
      6'b100001 : _zz_shift_q_6_4 = shift_q_map_33;
      6'b100010 : _zz_shift_q_6_4 = shift_q_map_34;
      6'b100011 : _zz_shift_q_6_4 = shift_q_map_35;
      6'b100100 : _zz_shift_q_6_4 = shift_q_map_36;
      6'b100101 : _zz_shift_q_6_4 = shift_q_map_37;
      6'b100110 : _zz_shift_q_6_4 = shift_q_map_38;
      6'b100111 : _zz_shift_q_6_4 = shift_q_map_39;
      6'b101000 : _zz_shift_q_6_4 = shift_q_map_40;
      6'b101001 : _zz_shift_q_6_4 = shift_q_map_41;
      6'b101010 : _zz_shift_q_6_4 = shift_q_map_42;
      6'b101011 : _zz_shift_q_6_4 = shift_q_map_43;
      6'b101100 : _zz_shift_q_6_4 = shift_q_map_44;
      6'b101101 : _zz_shift_q_6_4 = shift_q_map_45;
      6'b101110 : _zz_shift_q_6_4 = shift_q_map_46;
      6'b101111 : _zz_shift_q_6_4 = shift_q_map_47;
      6'b110000 : _zz_shift_q_6_4 = shift_q_map_48;
      6'b110001 : _zz_shift_q_6_4 = shift_q_map_49;
      6'b110010 : _zz_shift_q_6_4 = shift_q_map_50;
      6'b110011 : _zz_shift_q_6_4 = shift_q_map_51;
      6'b110100 : _zz_shift_q_6_4 = shift_q_map_52;
      6'b110101 : _zz_shift_q_6_4 = shift_q_map_53;
      6'b110110 : _zz_shift_q_6_4 = shift_q_map_54;
      6'b110111 : _zz_shift_q_6_4 = shift_q_map_55;
      6'b111000 : _zz_shift_q_6_4 = shift_q_map_56;
      6'b111001 : _zz_shift_q_6_4 = shift_q_map_57;
      6'b111010 : _zz_shift_q_6_4 = shift_q_map_58;
      6'b111011 : _zz_shift_q_6_4 = shift_q_map_59;
      6'b111100 : _zz_shift_q_6_4 = shift_q_map_60;
      6'b111101 : _zz_shift_q_6_4 = shift_q_map_61;
      6'b111110 : _zz_shift_q_6_4 = shift_q_map_62;
      default : _zz_shift_q_6_4 = shift_q_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_7_5)
      6'b000000 : _zz_shift_i_7_4 = shift_i_map_0;
      6'b000001 : _zz_shift_i_7_4 = shift_i_map_1;
      6'b000010 : _zz_shift_i_7_4 = shift_i_map_2;
      6'b000011 : _zz_shift_i_7_4 = shift_i_map_3;
      6'b000100 : _zz_shift_i_7_4 = shift_i_map_4;
      6'b000101 : _zz_shift_i_7_4 = shift_i_map_5;
      6'b000110 : _zz_shift_i_7_4 = shift_i_map_6;
      6'b000111 : _zz_shift_i_7_4 = shift_i_map_7;
      6'b001000 : _zz_shift_i_7_4 = shift_i_map_8;
      6'b001001 : _zz_shift_i_7_4 = shift_i_map_9;
      6'b001010 : _zz_shift_i_7_4 = shift_i_map_10;
      6'b001011 : _zz_shift_i_7_4 = shift_i_map_11;
      6'b001100 : _zz_shift_i_7_4 = shift_i_map_12;
      6'b001101 : _zz_shift_i_7_4 = shift_i_map_13;
      6'b001110 : _zz_shift_i_7_4 = shift_i_map_14;
      6'b001111 : _zz_shift_i_7_4 = shift_i_map_15;
      6'b010000 : _zz_shift_i_7_4 = shift_i_map_16;
      6'b010001 : _zz_shift_i_7_4 = shift_i_map_17;
      6'b010010 : _zz_shift_i_7_4 = shift_i_map_18;
      6'b010011 : _zz_shift_i_7_4 = shift_i_map_19;
      6'b010100 : _zz_shift_i_7_4 = shift_i_map_20;
      6'b010101 : _zz_shift_i_7_4 = shift_i_map_21;
      6'b010110 : _zz_shift_i_7_4 = shift_i_map_22;
      6'b010111 : _zz_shift_i_7_4 = shift_i_map_23;
      6'b011000 : _zz_shift_i_7_4 = shift_i_map_24;
      6'b011001 : _zz_shift_i_7_4 = shift_i_map_25;
      6'b011010 : _zz_shift_i_7_4 = shift_i_map_26;
      6'b011011 : _zz_shift_i_7_4 = shift_i_map_27;
      6'b011100 : _zz_shift_i_7_4 = shift_i_map_28;
      6'b011101 : _zz_shift_i_7_4 = shift_i_map_29;
      6'b011110 : _zz_shift_i_7_4 = shift_i_map_30;
      6'b011111 : _zz_shift_i_7_4 = shift_i_map_31;
      6'b100000 : _zz_shift_i_7_4 = shift_i_map_32;
      6'b100001 : _zz_shift_i_7_4 = shift_i_map_33;
      6'b100010 : _zz_shift_i_7_4 = shift_i_map_34;
      6'b100011 : _zz_shift_i_7_4 = shift_i_map_35;
      6'b100100 : _zz_shift_i_7_4 = shift_i_map_36;
      6'b100101 : _zz_shift_i_7_4 = shift_i_map_37;
      6'b100110 : _zz_shift_i_7_4 = shift_i_map_38;
      6'b100111 : _zz_shift_i_7_4 = shift_i_map_39;
      6'b101000 : _zz_shift_i_7_4 = shift_i_map_40;
      6'b101001 : _zz_shift_i_7_4 = shift_i_map_41;
      6'b101010 : _zz_shift_i_7_4 = shift_i_map_42;
      6'b101011 : _zz_shift_i_7_4 = shift_i_map_43;
      6'b101100 : _zz_shift_i_7_4 = shift_i_map_44;
      6'b101101 : _zz_shift_i_7_4 = shift_i_map_45;
      6'b101110 : _zz_shift_i_7_4 = shift_i_map_46;
      6'b101111 : _zz_shift_i_7_4 = shift_i_map_47;
      6'b110000 : _zz_shift_i_7_4 = shift_i_map_48;
      6'b110001 : _zz_shift_i_7_4 = shift_i_map_49;
      6'b110010 : _zz_shift_i_7_4 = shift_i_map_50;
      6'b110011 : _zz_shift_i_7_4 = shift_i_map_51;
      6'b110100 : _zz_shift_i_7_4 = shift_i_map_52;
      6'b110101 : _zz_shift_i_7_4 = shift_i_map_53;
      6'b110110 : _zz_shift_i_7_4 = shift_i_map_54;
      6'b110111 : _zz_shift_i_7_4 = shift_i_map_55;
      6'b111000 : _zz_shift_i_7_4 = shift_i_map_56;
      6'b111001 : _zz_shift_i_7_4 = shift_i_map_57;
      6'b111010 : _zz_shift_i_7_4 = shift_i_map_58;
      6'b111011 : _zz_shift_i_7_4 = shift_i_map_59;
      6'b111100 : _zz_shift_i_7_4 = shift_i_map_60;
      6'b111101 : _zz_shift_i_7_4 = shift_i_map_61;
      6'b111110 : _zz_shift_i_7_4 = shift_i_map_62;
      default : _zz_shift_i_7_4 = shift_i_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_7_5)
      6'b000000 : _zz_shift_q_7_4 = shift_q_map_0;
      6'b000001 : _zz_shift_q_7_4 = shift_q_map_1;
      6'b000010 : _zz_shift_q_7_4 = shift_q_map_2;
      6'b000011 : _zz_shift_q_7_4 = shift_q_map_3;
      6'b000100 : _zz_shift_q_7_4 = shift_q_map_4;
      6'b000101 : _zz_shift_q_7_4 = shift_q_map_5;
      6'b000110 : _zz_shift_q_7_4 = shift_q_map_6;
      6'b000111 : _zz_shift_q_7_4 = shift_q_map_7;
      6'b001000 : _zz_shift_q_7_4 = shift_q_map_8;
      6'b001001 : _zz_shift_q_7_4 = shift_q_map_9;
      6'b001010 : _zz_shift_q_7_4 = shift_q_map_10;
      6'b001011 : _zz_shift_q_7_4 = shift_q_map_11;
      6'b001100 : _zz_shift_q_7_4 = shift_q_map_12;
      6'b001101 : _zz_shift_q_7_4 = shift_q_map_13;
      6'b001110 : _zz_shift_q_7_4 = shift_q_map_14;
      6'b001111 : _zz_shift_q_7_4 = shift_q_map_15;
      6'b010000 : _zz_shift_q_7_4 = shift_q_map_16;
      6'b010001 : _zz_shift_q_7_4 = shift_q_map_17;
      6'b010010 : _zz_shift_q_7_4 = shift_q_map_18;
      6'b010011 : _zz_shift_q_7_4 = shift_q_map_19;
      6'b010100 : _zz_shift_q_7_4 = shift_q_map_20;
      6'b010101 : _zz_shift_q_7_4 = shift_q_map_21;
      6'b010110 : _zz_shift_q_7_4 = shift_q_map_22;
      6'b010111 : _zz_shift_q_7_4 = shift_q_map_23;
      6'b011000 : _zz_shift_q_7_4 = shift_q_map_24;
      6'b011001 : _zz_shift_q_7_4 = shift_q_map_25;
      6'b011010 : _zz_shift_q_7_4 = shift_q_map_26;
      6'b011011 : _zz_shift_q_7_4 = shift_q_map_27;
      6'b011100 : _zz_shift_q_7_4 = shift_q_map_28;
      6'b011101 : _zz_shift_q_7_4 = shift_q_map_29;
      6'b011110 : _zz_shift_q_7_4 = shift_q_map_30;
      6'b011111 : _zz_shift_q_7_4 = shift_q_map_31;
      6'b100000 : _zz_shift_q_7_4 = shift_q_map_32;
      6'b100001 : _zz_shift_q_7_4 = shift_q_map_33;
      6'b100010 : _zz_shift_q_7_4 = shift_q_map_34;
      6'b100011 : _zz_shift_q_7_4 = shift_q_map_35;
      6'b100100 : _zz_shift_q_7_4 = shift_q_map_36;
      6'b100101 : _zz_shift_q_7_4 = shift_q_map_37;
      6'b100110 : _zz_shift_q_7_4 = shift_q_map_38;
      6'b100111 : _zz_shift_q_7_4 = shift_q_map_39;
      6'b101000 : _zz_shift_q_7_4 = shift_q_map_40;
      6'b101001 : _zz_shift_q_7_4 = shift_q_map_41;
      6'b101010 : _zz_shift_q_7_4 = shift_q_map_42;
      6'b101011 : _zz_shift_q_7_4 = shift_q_map_43;
      6'b101100 : _zz_shift_q_7_4 = shift_q_map_44;
      6'b101101 : _zz_shift_q_7_4 = shift_q_map_45;
      6'b101110 : _zz_shift_q_7_4 = shift_q_map_46;
      6'b101111 : _zz_shift_q_7_4 = shift_q_map_47;
      6'b110000 : _zz_shift_q_7_4 = shift_q_map_48;
      6'b110001 : _zz_shift_q_7_4 = shift_q_map_49;
      6'b110010 : _zz_shift_q_7_4 = shift_q_map_50;
      6'b110011 : _zz_shift_q_7_4 = shift_q_map_51;
      6'b110100 : _zz_shift_q_7_4 = shift_q_map_52;
      6'b110101 : _zz_shift_q_7_4 = shift_q_map_53;
      6'b110110 : _zz_shift_q_7_4 = shift_q_map_54;
      6'b110111 : _zz_shift_q_7_4 = shift_q_map_55;
      6'b111000 : _zz_shift_q_7_4 = shift_q_map_56;
      6'b111001 : _zz_shift_q_7_4 = shift_q_map_57;
      6'b111010 : _zz_shift_q_7_4 = shift_q_map_58;
      6'b111011 : _zz_shift_q_7_4 = shift_q_map_59;
      6'b111100 : _zz_shift_q_7_4 = shift_q_map_60;
      6'b111101 : _zz_shift_q_7_4 = shift_q_map_61;
      6'b111110 : _zz_shift_q_7_4 = shift_q_map_62;
      default : _zz_shift_q_7_4 = shift_q_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_0_7)
      6'b000000 : _zz_shift_i_0_6 = shift_i_map_0;
      6'b000001 : _zz_shift_i_0_6 = shift_i_map_1;
      6'b000010 : _zz_shift_i_0_6 = shift_i_map_2;
      6'b000011 : _zz_shift_i_0_6 = shift_i_map_3;
      6'b000100 : _zz_shift_i_0_6 = shift_i_map_4;
      6'b000101 : _zz_shift_i_0_6 = shift_i_map_5;
      6'b000110 : _zz_shift_i_0_6 = shift_i_map_6;
      6'b000111 : _zz_shift_i_0_6 = shift_i_map_7;
      6'b001000 : _zz_shift_i_0_6 = shift_i_map_8;
      6'b001001 : _zz_shift_i_0_6 = shift_i_map_9;
      6'b001010 : _zz_shift_i_0_6 = shift_i_map_10;
      6'b001011 : _zz_shift_i_0_6 = shift_i_map_11;
      6'b001100 : _zz_shift_i_0_6 = shift_i_map_12;
      6'b001101 : _zz_shift_i_0_6 = shift_i_map_13;
      6'b001110 : _zz_shift_i_0_6 = shift_i_map_14;
      6'b001111 : _zz_shift_i_0_6 = shift_i_map_15;
      6'b010000 : _zz_shift_i_0_6 = shift_i_map_16;
      6'b010001 : _zz_shift_i_0_6 = shift_i_map_17;
      6'b010010 : _zz_shift_i_0_6 = shift_i_map_18;
      6'b010011 : _zz_shift_i_0_6 = shift_i_map_19;
      6'b010100 : _zz_shift_i_0_6 = shift_i_map_20;
      6'b010101 : _zz_shift_i_0_6 = shift_i_map_21;
      6'b010110 : _zz_shift_i_0_6 = shift_i_map_22;
      6'b010111 : _zz_shift_i_0_6 = shift_i_map_23;
      6'b011000 : _zz_shift_i_0_6 = shift_i_map_24;
      6'b011001 : _zz_shift_i_0_6 = shift_i_map_25;
      6'b011010 : _zz_shift_i_0_6 = shift_i_map_26;
      6'b011011 : _zz_shift_i_0_6 = shift_i_map_27;
      6'b011100 : _zz_shift_i_0_6 = shift_i_map_28;
      6'b011101 : _zz_shift_i_0_6 = shift_i_map_29;
      6'b011110 : _zz_shift_i_0_6 = shift_i_map_30;
      6'b011111 : _zz_shift_i_0_6 = shift_i_map_31;
      6'b100000 : _zz_shift_i_0_6 = shift_i_map_32;
      6'b100001 : _zz_shift_i_0_6 = shift_i_map_33;
      6'b100010 : _zz_shift_i_0_6 = shift_i_map_34;
      6'b100011 : _zz_shift_i_0_6 = shift_i_map_35;
      6'b100100 : _zz_shift_i_0_6 = shift_i_map_36;
      6'b100101 : _zz_shift_i_0_6 = shift_i_map_37;
      6'b100110 : _zz_shift_i_0_6 = shift_i_map_38;
      6'b100111 : _zz_shift_i_0_6 = shift_i_map_39;
      6'b101000 : _zz_shift_i_0_6 = shift_i_map_40;
      6'b101001 : _zz_shift_i_0_6 = shift_i_map_41;
      6'b101010 : _zz_shift_i_0_6 = shift_i_map_42;
      6'b101011 : _zz_shift_i_0_6 = shift_i_map_43;
      6'b101100 : _zz_shift_i_0_6 = shift_i_map_44;
      6'b101101 : _zz_shift_i_0_6 = shift_i_map_45;
      6'b101110 : _zz_shift_i_0_6 = shift_i_map_46;
      6'b101111 : _zz_shift_i_0_6 = shift_i_map_47;
      6'b110000 : _zz_shift_i_0_6 = shift_i_map_48;
      6'b110001 : _zz_shift_i_0_6 = shift_i_map_49;
      6'b110010 : _zz_shift_i_0_6 = shift_i_map_50;
      6'b110011 : _zz_shift_i_0_6 = shift_i_map_51;
      6'b110100 : _zz_shift_i_0_6 = shift_i_map_52;
      6'b110101 : _zz_shift_i_0_6 = shift_i_map_53;
      6'b110110 : _zz_shift_i_0_6 = shift_i_map_54;
      6'b110111 : _zz_shift_i_0_6 = shift_i_map_55;
      6'b111000 : _zz_shift_i_0_6 = shift_i_map_56;
      6'b111001 : _zz_shift_i_0_6 = shift_i_map_57;
      6'b111010 : _zz_shift_i_0_6 = shift_i_map_58;
      6'b111011 : _zz_shift_i_0_6 = shift_i_map_59;
      6'b111100 : _zz_shift_i_0_6 = shift_i_map_60;
      6'b111101 : _zz_shift_i_0_6 = shift_i_map_61;
      6'b111110 : _zz_shift_i_0_6 = shift_i_map_62;
      default : _zz_shift_i_0_6 = shift_i_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_0_7)
      6'b000000 : _zz_shift_q_0_6 = shift_q_map_0;
      6'b000001 : _zz_shift_q_0_6 = shift_q_map_1;
      6'b000010 : _zz_shift_q_0_6 = shift_q_map_2;
      6'b000011 : _zz_shift_q_0_6 = shift_q_map_3;
      6'b000100 : _zz_shift_q_0_6 = shift_q_map_4;
      6'b000101 : _zz_shift_q_0_6 = shift_q_map_5;
      6'b000110 : _zz_shift_q_0_6 = shift_q_map_6;
      6'b000111 : _zz_shift_q_0_6 = shift_q_map_7;
      6'b001000 : _zz_shift_q_0_6 = shift_q_map_8;
      6'b001001 : _zz_shift_q_0_6 = shift_q_map_9;
      6'b001010 : _zz_shift_q_0_6 = shift_q_map_10;
      6'b001011 : _zz_shift_q_0_6 = shift_q_map_11;
      6'b001100 : _zz_shift_q_0_6 = shift_q_map_12;
      6'b001101 : _zz_shift_q_0_6 = shift_q_map_13;
      6'b001110 : _zz_shift_q_0_6 = shift_q_map_14;
      6'b001111 : _zz_shift_q_0_6 = shift_q_map_15;
      6'b010000 : _zz_shift_q_0_6 = shift_q_map_16;
      6'b010001 : _zz_shift_q_0_6 = shift_q_map_17;
      6'b010010 : _zz_shift_q_0_6 = shift_q_map_18;
      6'b010011 : _zz_shift_q_0_6 = shift_q_map_19;
      6'b010100 : _zz_shift_q_0_6 = shift_q_map_20;
      6'b010101 : _zz_shift_q_0_6 = shift_q_map_21;
      6'b010110 : _zz_shift_q_0_6 = shift_q_map_22;
      6'b010111 : _zz_shift_q_0_6 = shift_q_map_23;
      6'b011000 : _zz_shift_q_0_6 = shift_q_map_24;
      6'b011001 : _zz_shift_q_0_6 = shift_q_map_25;
      6'b011010 : _zz_shift_q_0_6 = shift_q_map_26;
      6'b011011 : _zz_shift_q_0_6 = shift_q_map_27;
      6'b011100 : _zz_shift_q_0_6 = shift_q_map_28;
      6'b011101 : _zz_shift_q_0_6 = shift_q_map_29;
      6'b011110 : _zz_shift_q_0_6 = shift_q_map_30;
      6'b011111 : _zz_shift_q_0_6 = shift_q_map_31;
      6'b100000 : _zz_shift_q_0_6 = shift_q_map_32;
      6'b100001 : _zz_shift_q_0_6 = shift_q_map_33;
      6'b100010 : _zz_shift_q_0_6 = shift_q_map_34;
      6'b100011 : _zz_shift_q_0_6 = shift_q_map_35;
      6'b100100 : _zz_shift_q_0_6 = shift_q_map_36;
      6'b100101 : _zz_shift_q_0_6 = shift_q_map_37;
      6'b100110 : _zz_shift_q_0_6 = shift_q_map_38;
      6'b100111 : _zz_shift_q_0_6 = shift_q_map_39;
      6'b101000 : _zz_shift_q_0_6 = shift_q_map_40;
      6'b101001 : _zz_shift_q_0_6 = shift_q_map_41;
      6'b101010 : _zz_shift_q_0_6 = shift_q_map_42;
      6'b101011 : _zz_shift_q_0_6 = shift_q_map_43;
      6'b101100 : _zz_shift_q_0_6 = shift_q_map_44;
      6'b101101 : _zz_shift_q_0_6 = shift_q_map_45;
      6'b101110 : _zz_shift_q_0_6 = shift_q_map_46;
      6'b101111 : _zz_shift_q_0_6 = shift_q_map_47;
      6'b110000 : _zz_shift_q_0_6 = shift_q_map_48;
      6'b110001 : _zz_shift_q_0_6 = shift_q_map_49;
      6'b110010 : _zz_shift_q_0_6 = shift_q_map_50;
      6'b110011 : _zz_shift_q_0_6 = shift_q_map_51;
      6'b110100 : _zz_shift_q_0_6 = shift_q_map_52;
      6'b110101 : _zz_shift_q_0_6 = shift_q_map_53;
      6'b110110 : _zz_shift_q_0_6 = shift_q_map_54;
      6'b110111 : _zz_shift_q_0_6 = shift_q_map_55;
      6'b111000 : _zz_shift_q_0_6 = shift_q_map_56;
      6'b111001 : _zz_shift_q_0_6 = shift_q_map_57;
      6'b111010 : _zz_shift_q_0_6 = shift_q_map_58;
      6'b111011 : _zz_shift_q_0_6 = shift_q_map_59;
      6'b111100 : _zz_shift_q_0_6 = shift_q_map_60;
      6'b111101 : _zz_shift_q_0_6 = shift_q_map_61;
      6'b111110 : _zz_shift_q_0_6 = shift_q_map_62;
      default : _zz_shift_q_0_6 = shift_q_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_1_7)
      6'b000000 : _zz_shift_i_1_6 = shift_i_map_0;
      6'b000001 : _zz_shift_i_1_6 = shift_i_map_1;
      6'b000010 : _zz_shift_i_1_6 = shift_i_map_2;
      6'b000011 : _zz_shift_i_1_6 = shift_i_map_3;
      6'b000100 : _zz_shift_i_1_6 = shift_i_map_4;
      6'b000101 : _zz_shift_i_1_6 = shift_i_map_5;
      6'b000110 : _zz_shift_i_1_6 = shift_i_map_6;
      6'b000111 : _zz_shift_i_1_6 = shift_i_map_7;
      6'b001000 : _zz_shift_i_1_6 = shift_i_map_8;
      6'b001001 : _zz_shift_i_1_6 = shift_i_map_9;
      6'b001010 : _zz_shift_i_1_6 = shift_i_map_10;
      6'b001011 : _zz_shift_i_1_6 = shift_i_map_11;
      6'b001100 : _zz_shift_i_1_6 = shift_i_map_12;
      6'b001101 : _zz_shift_i_1_6 = shift_i_map_13;
      6'b001110 : _zz_shift_i_1_6 = shift_i_map_14;
      6'b001111 : _zz_shift_i_1_6 = shift_i_map_15;
      6'b010000 : _zz_shift_i_1_6 = shift_i_map_16;
      6'b010001 : _zz_shift_i_1_6 = shift_i_map_17;
      6'b010010 : _zz_shift_i_1_6 = shift_i_map_18;
      6'b010011 : _zz_shift_i_1_6 = shift_i_map_19;
      6'b010100 : _zz_shift_i_1_6 = shift_i_map_20;
      6'b010101 : _zz_shift_i_1_6 = shift_i_map_21;
      6'b010110 : _zz_shift_i_1_6 = shift_i_map_22;
      6'b010111 : _zz_shift_i_1_6 = shift_i_map_23;
      6'b011000 : _zz_shift_i_1_6 = shift_i_map_24;
      6'b011001 : _zz_shift_i_1_6 = shift_i_map_25;
      6'b011010 : _zz_shift_i_1_6 = shift_i_map_26;
      6'b011011 : _zz_shift_i_1_6 = shift_i_map_27;
      6'b011100 : _zz_shift_i_1_6 = shift_i_map_28;
      6'b011101 : _zz_shift_i_1_6 = shift_i_map_29;
      6'b011110 : _zz_shift_i_1_6 = shift_i_map_30;
      6'b011111 : _zz_shift_i_1_6 = shift_i_map_31;
      6'b100000 : _zz_shift_i_1_6 = shift_i_map_32;
      6'b100001 : _zz_shift_i_1_6 = shift_i_map_33;
      6'b100010 : _zz_shift_i_1_6 = shift_i_map_34;
      6'b100011 : _zz_shift_i_1_6 = shift_i_map_35;
      6'b100100 : _zz_shift_i_1_6 = shift_i_map_36;
      6'b100101 : _zz_shift_i_1_6 = shift_i_map_37;
      6'b100110 : _zz_shift_i_1_6 = shift_i_map_38;
      6'b100111 : _zz_shift_i_1_6 = shift_i_map_39;
      6'b101000 : _zz_shift_i_1_6 = shift_i_map_40;
      6'b101001 : _zz_shift_i_1_6 = shift_i_map_41;
      6'b101010 : _zz_shift_i_1_6 = shift_i_map_42;
      6'b101011 : _zz_shift_i_1_6 = shift_i_map_43;
      6'b101100 : _zz_shift_i_1_6 = shift_i_map_44;
      6'b101101 : _zz_shift_i_1_6 = shift_i_map_45;
      6'b101110 : _zz_shift_i_1_6 = shift_i_map_46;
      6'b101111 : _zz_shift_i_1_6 = shift_i_map_47;
      6'b110000 : _zz_shift_i_1_6 = shift_i_map_48;
      6'b110001 : _zz_shift_i_1_6 = shift_i_map_49;
      6'b110010 : _zz_shift_i_1_6 = shift_i_map_50;
      6'b110011 : _zz_shift_i_1_6 = shift_i_map_51;
      6'b110100 : _zz_shift_i_1_6 = shift_i_map_52;
      6'b110101 : _zz_shift_i_1_6 = shift_i_map_53;
      6'b110110 : _zz_shift_i_1_6 = shift_i_map_54;
      6'b110111 : _zz_shift_i_1_6 = shift_i_map_55;
      6'b111000 : _zz_shift_i_1_6 = shift_i_map_56;
      6'b111001 : _zz_shift_i_1_6 = shift_i_map_57;
      6'b111010 : _zz_shift_i_1_6 = shift_i_map_58;
      6'b111011 : _zz_shift_i_1_6 = shift_i_map_59;
      6'b111100 : _zz_shift_i_1_6 = shift_i_map_60;
      6'b111101 : _zz_shift_i_1_6 = shift_i_map_61;
      6'b111110 : _zz_shift_i_1_6 = shift_i_map_62;
      default : _zz_shift_i_1_6 = shift_i_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_1_7)
      6'b000000 : _zz_shift_q_1_6 = shift_q_map_0;
      6'b000001 : _zz_shift_q_1_6 = shift_q_map_1;
      6'b000010 : _zz_shift_q_1_6 = shift_q_map_2;
      6'b000011 : _zz_shift_q_1_6 = shift_q_map_3;
      6'b000100 : _zz_shift_q_1_6 = shift_q_map_4;
      6'b000101 : _zz_shift_q_1_6 = shift_q_map_5;
      6'b000110 : _zz_shift_q_1_6 = shift_q_map_6;
      6'b000111 : _zz_shift_q_1_6 = shift_q_map_7;
      6'b001000 : _zz_shift_q_1_6 = shift_q_map_8;
      6'b001001 : _zz_shift_q_1_6 = shift_q_map_9;
      6'b001010 : _zz_shift_q_1_6 = shift_q_map_10;
      6'b001011 : _zz_shift_q_1_6 = shift_q_map_11;
      6'b001100 : _zz_shift_q_1_6 = shift_q_map_12;
      6'b001101 : _zz_shift_q_1_6 = shift_q_map_13;
      6'b001110 : _zz_shift_q_1_6 = shift_q_map_14;
      6'b001111 : _zz_shift_q_1_6 = shift_q_map_15;
      6'b010000 : _zz_shift_q_1_6 = shift_q_map_16;
      6'b010001 : _zz_shift_q_1_6 = shift_q_map_17;
      6'b010010 : _zz_shift_q_1_6 = shift_q_map_18;
      6'b010011 : _zz_shift_q_1_6 = shift_q_map_19;
      6'b010100 : _zz_shift_q_1_6 = shift_q_map_20;
      6'b010101 : _zz_shift_q_1_6 = shift_q_map_21;
      6'b010110 : _zz_shift_q_1_6 = shift_q_map_22;
      6'b010111 : _zz_shift_q_1_6 = shift_q_map_23;
      6'b011000 : _zz_shift_q_1_6 = shift_q_map_24;
      6'b011001 : _zz_shift_q_1_6 = shift_q_map_25;
      6'b011010 : _zz_shift_q_1_6 = shift_q_map_26;
      6'b011011 : _zz_shift_q_1_6 = shift_q_map_27;
      6'b011100 : _zz_shift_q_1_6 = shift_q_map_28;
      6'b011101 : _zz_shift_q_1_6 = shift_q_map_29;
      6'b011110 : _zz_shift_q_1_6 = shift_q_map_30;
      6'b011111 : _zz_shift_q_1_6 = shift_q_map_31;
      6'b100000 : _zz_shift_q_1_6 = shift_q_map_32;
      6'b100001 : _zz_shift_q_1_6 = shift_q_map_33;
      6'b100010 : _zz_shift_q_1_6 = shift_q_map_34;
      6'b100011 : _zz_shift_q_1_6 = shift_q_map_35;
      6'b100100 : _zz_shift_q_1_6 = shift_q_map_36;
      6'b100101 : _zz_shift_q_1_6 = shift_q_map_37;
      6'b100110 : _zz_shift_q_1_6 = shift_q_map_38;
      6'b100111 : _zz_shift_q_1_6 = shift_q_map_39;
      6'b101000 : _zz_shift_q_1_6 = shift_q_map_40;
      6'b101001 : _zz_shift_q_1_6 = shift_q_map_41;
      6'b101010 : _zz_shift_q_1_6 = shift_q_map_42;
      6'b101011 : _zz_shift_q_1_6 = shift_q_map_43;
      6'b101100 : _zz_shift_q_1_6 = shift_q_map_44;
      6'b101101 : _zz_shift_q_1_6 = shift_q_map_45;
      6'b101110 : _zz_shift_q_1_6 = shift_q_map_46;
      6'b101111 : _zz_shift_q_1_6 = shift_q_map_47;
      6'b110000 : _zz_shift_q_1_6 = shift_q_map_48;
      6'b110001 : _zz_shift_q_1_6 = shift_q_map_49;
      6'b110010 : _zz_shift_q_1_6 = shift_q_map_50;
      6'b110011 : _zz_shift_q_1_6 = shift_q_map_51;
      6'b110100 : _zz_shift_q_1_6 = shift_q_map_52;
      6'b110101 : _zz_shift_q_1_6 = shift_q_map_53;
      6'b110110 : _zz_shift_q_1_6 = shift_q_map_54;
      6'b110111 : _zz_shift_q_1_6 = shift_q_map_55;
      6'b111000 : _zz_shift_q_1_6 = shift_q_map_56;
      6'b111001 : _zz_shift_q_1_6 = shift_q_map_57;
      6'b111010 : _zz_shift_q_1_6 = shift_q_map_58;
      6'b111011 : _zz_shift_q_1_6 = shift_q_map_59;
      6'b111100 : _zz_shift_q_1_6 = shift_q_map_60;
      6'b111101 : _zz_shift_q_1_6 = shift_q_map_61;
      6'b111110 : _zz_shift_q_1_6 = shift_q_map_62;
      default : _zz_shift_q_1_6 = shift_q_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_2_7)
      6'b000000 : _zz_shift_i_2_6 = shift_i_map_0;
      6'b000001 : _zz_shift_i_2_6 = shift_i_map_1;
      6'b000010 : _zz_shift_i_2_6 = shift_i_map_2;
      6'b000011 : _zz_shift_i_2_6 = shift_i_map_3;
      6'b000100 : _zz_shift_i_2_6 = shift_i_map_4;
      6'b000101 : _zz_shift_i_2_6 = shift_i_map_5;
      6'b000110 : _zz_shift_i_2_6 = shift_i_map_6;
      6'b000111 : _zz_shift_i_2_6 = shift_i_map_7;
      6'b001000 : _zz_shift_i_2_6 = shift_i_map_8;
      6'b001001 : _zz_shift_i_2_6 = shift_i_map_9;
      6'b001010 : _zz_shift_i_2_6 = shift_i_map_10;
      6'b001011 : _zz_shift_i_2_6 = shift_i_map_11;
      6'b001100 : _zz_shift_i_2_6 = shift_i_map_12;
      6'b001101 : _zz_shift_i_2_6 = shift_i_map_13;
      6'b001110 : _zz_shift_i_2_6 = shift_i_map_14;
      6'b001111 : _zz_shift_i_2_6 = shift_i_map_15;
      6'b010000 : _zz_shift_i_2_6 = shift_i_map_16;
      6'b010001 : _zz_shift_i_2_6 = shift_i_map_17;
      6'b010010 : _zz_shift_i_2_6 = shift_i_map_18;
      6'b010011 : _zz_shift_i_2_6 = shift_i_map_19;
      6'b010100 : _zz_shift_i_2_6 = shift_i_map_20;
      6'b010101 : _zz_shift_i_2_6 = shift_i_map_21;
      6'b010110 : _zz_shift_i_2_6 = shift_i_map_22;
      6'b010111 : _zz_shift_i_2_6 = shift_i_map_23;
      6'b011000 : _zz_shift_i_2_6 = shift_i_map_24;
      6'b011001 : _zz_shift_i_2_6 = shift_i_map_25;
      6'b011010 : _zz_shift_i_2_6 = shift_i_map_26;
      6'b011011 : _zz_shift_i_2_6 = shift_i_map_27;
      6'b011100 : _zz_shift_i_2_6 = shift_i_map_28;
      6'b011101 : _zz_shift_i_2_6 = shift_i_map_29;
      6'b011110 : _zz_shift_i_2_6 = shift_i_map_30;
      6'b011111 : _zz_shift_i_2_6 = shift_i_map_31;
      6'b100000 : _zz_shift_i_2_6 = shift_i_map_32;
      6'b100001 : _zz_shift_i_2_6 = shift_i_map_33;
      6'b100010 : _zz_shift_i_2_6 = shift_i_map_34;
      6'b100011 : _zz_shift_i_2_6 = shift_i_map_35;
      6'b100100 : _zz_shift_i_2_6 = shift_i_map_36;
      6'b100101 : _zz_shift_i_2_6 = shift_i_map_37;
      6'b100110 : _zz_shift_i_2_6 = shift_i_map_38;
      6'b100111 : _zz_shift_i_2_6 = shift_i_map_39;
      6'b101000 : _zz_shift_i_2_6 = shift_i_map_40;
      6'b101001 : _zz_shift_i_2_6 = shift_i_map_41;
      6'b101010 : _zz_shift_i_2_6 = shift_i_map_42;
      6'b101011 : _zz_shift_i_2_6 = shift_i_map_43;
      6'b101100 : _zz_shift_i_2_6 = shift_i_map_44;
      6'b101101 : _zz_shift_i_2_6 = shift_i_map_45;
      6'b101110 : _zz_shift_i_2_6 = shift_i_map_46;
      6'b101111 : _zz_shift_i_2_6 = shift_i_map_47;
      6'b110000 : _zz_shift_i_2_6 = shift_i_map_48;
      6'b110001 : _zz_shift_i_2_6 = shift_i_map_49;
      6'b110010 : _zz_shift_i_2_6 = shift_i_map_50;
      6'b110011 : _zz_shift_i_2_6 = shift_i_map_51;
      6'b110100 : _zz_shift_i_2_6 = shift_i_map_52;
      6'b110101 : _zz_shift_i_2_6 = shift_i_map_53;
      6'b110110 : _zz_shift_i_2_6 = shift_i_map_54;
      6'b110111 : _zz_shift_i_2_6 = shift_i_map_55;
      6'b111000 : _zz_shift_i_2_6 = shift_i_map_56;
      6'b111001 : _zz_shift_i_2_6 = shift_i_map_57;
      6'b111010 : _zz_shift_i_2_6 = shift_i_map_58;
      6'b111011 : _zz_shift_i_2_6 = shift_i_map_59;
      6'b111100 : _zz_shift_i_2_6 = shift_i_map_60;
      6'b111101 : _zz_shift_i_2_6 = shift_i_map_61;
      6'b111110 : _zz_shift_i_2_6 = shift_i_map_62;
      default : _zz_shift_i_2_6 = shift_i_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_2_7)
      6'b000000 : _zz_shift_q_2_6 = shift_q_map_0;
      6'b000001 : _zz_shift_q_2_6 = shift_q_map_1;
      6'b000010 : _zz_shift_q_2_6 = shift_q_map_2;
      6'b000011 : _zz_shift_q_2_6 = shift_q_map_3;
      6'b000100 : _zz_shift_q_2_6 = shift_q_map_4;
      6'b000101 : _zz_shift_q_2_6 = shift_q_map_5;
      6'b000110 : _zz_shift_q_2_6 = shift_q_map_6;
      6'b000111 : _zz_shift_q_2_6 = shift_q_map_7;
      6'b001000 : _zz_shift_q_2_6 = shift_q_map_8;
      6'b001001 : _zz_shift_q_2_6 = shift_q_map_9;
      6'b001010 : _zz_shift_q_2_6 = shift_q_map_10;
      6'b001011 : _zz_shift_q_2_6 = shift_q_map_11;
      6'b001100 : _zz_shift_q_2_6 = shift_q_map_12;
      6'b001101 : _zz_shift_q_2_6 = shift_q_map_13;
      6'b001110 : _zz_shift_q_2_6 = shift_q_map_14;
      6'b001111 : _zz_shift_q_2_6 = shift_q_map_15;
      6'b010000 : _zz_shift_q_2_6 = shift_q_map_16;
      6'b010001 : _zz_shift_q_2_6 = shift_q_map_17;
      6'b010010 : _zz_shift_q_2_6 = shift_q_map_18;
      6'b010011 : _zz_shift_q_2_6 = shift_q_map_19;
      6'b010100 : _zz_shift_q_2_6 = shift_q_map_20;
      6'b010101 : _zz_shift_q_2_6 = shift_q_map_21;
      6'b010110 : _zz_shift_q_2_6 = shift_q_map_22;
      6'b010111 : _zz_shift_q_2_6 = shift_q_map_23;
      6'b011000 : _zz_shift_q_2_6 = shift_q_map_24;
      6'b011001 : _zz_shift_q_2_6 = shift_q_map_25;
      6'b011010 : _zz_shift_q_2_6 = shift_q_map_26;
      6'b011011 : _zz_shift_q_2_6 = shift_q_map_27;
      6'b011100 : _zz_shift_q_2_6 = shift_q_map_28;
      6'b011101 : _zz_shift_q_2_6 = shift_q_map_29;
      6'b011110 : _zz_shift_q_2_6 = shift_q_map_30;
      6'b011111 : _zz_shift_q_2_6 = shift_q_map_31;
      6'b100000 : _zz_shift_q_2_6 = shift_q_map_32;
      6'b100001 : _zz_shift_q_2_6 = shift_q_map_33;
      6'b100010 : _zz_shift_q_2_6 = shift_q_map_34;
      6'b100011 : _zz_shift_q_2_6 = shift_q_map_35;
      6'b100100 : _zz_shift_q_2_6 = shift_q_map_36;
      6'b100101 : _zz_shift_q_2_6 = shift_q_map_37;
      6'b100110 : _zz_shift_q_2_6 = shift_q_map_38;
      6'b100111 : _zz_shift_q_2_6 = shift_q_map_39;
      6'b101000 : _zz_shift_q_2_6 = shift_q_map_40;
      6'b101001 : _zz_shift_q_2_6 = shift_q_map_41;
      6'b101010 : _zz_shift_q_2_6 = shift_q_map_42;
      6'b101011 : _zz_shift_q_2_6 = shift_q_map_43;
      6'b101100 : _zz_shift_q_2_6 = shift_q_map_44;
      6'b101101 : _zz_shift_q_2_6 = shift_q_map_45;
      6'b101110 : _zz_shift_q_2_6 = shift_q_map_46;
      6'b101111 : _zz_shift_q_2_6 = shift_q_map_47;
      6'b110000 : _zz_shift_q_2_6 = shift_q_map_48;
      6'b110001 : _zz_shift_q_2_6 = shift_q_map_49;
      6'b110010 : _zz_shift_q_2_6 = shift_q_map_50;
      6'b110011 : _zz_shift_q_2_6 = shift_q_map_51;
      6'b110100 : _zz_shift_q_2_6 = shift_q_map_52;
      6'b110101 : _zz_shift_q_2_6 = shift_q_map_53;
      6'b110110 : _zz_shift_q_2_6 = shift_q_map_54;
      6'b110111 : _zz_shift_q_2_6 = shift_q_map_55;
      6'b111000 : _zz_shift_q_2_6 = shift_q_map_56;
      6'b111001 : _zz_shift_q_2_6 = shift_q_map_57;
      6'b111010 : _zz_shift_q_2_6 = shift_q_map_58;
      6'b111011 : _zz_shift_q_2_6 = shift_q_map_59;
      6'b111100 : _zz_shift_q_2_6 = shift_q_map_60;
      6'b111101 : _zz_shift_q_2_6 = shift_q_map_61;
      6'b111110 : _zz_shift_q_2_6 = shift_q_map_62;
      default : _zz_shift_q_2_6 = shift_q_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_3_7)
      6'b000000 : _zz_shift_i_3_6 = shift_i_map_0;
      6'b000001 : _zz_shift_i_3_6 = shift_i_map_1;
      6'b000010 : _zz_shift_i_3_6 = shift_i_map_2;
      6'b000011 : _zz_shift_i_3_6 = shift_i_map_3;
      6'b000100 : _zz_shift_i_3_6 = shift_i_map_4;
      6'b000101 : _zz_shift_i_3_6 = shift_i_map_5;
      6'b000110 : _zz_shift_i_3_6 = shift_i_map_6;
      6'b000111 : _zz_shift_i_3_6 = shift_i_map_7;
      6'b001000 : _zz_shift_i_3_6 = shift_i_map_8;
      6'b001001 : _zz_shift_i_3_6 = shift_i_map_9;
      6'b001010 : _zz_shift_i_3_6 = shift_i_map_10;
      6'b001011 : _zz_shift_i_3_6 = shift_i_map_11;
      6'b001100 : _zz_shift_i_3_6 = shift_i_map_12;
      6'b001101 : _zz_shift_i_3_6 = shift_i_map_13;
      6'b001110 : _zz_shift_i_3_6 = shift_i_map_14;
      6'b001111 : _zz_shift_i_3_6 = shift_i_map_15;
      6'b010000 : _zz_shift_i_3_6 = shift_i_map_16;
      6'b010001 : _zz_shift_i_3_6 = shift_i_map_17;
      6'b010010 : _zz_shift_i_3_6 = shift_i_map_18;
      6'b010011 : _zz_shift_i_3_6 = shift_i_map_19;
      6'b010100 : _zz_shift_i_3_6 = shift_i_map_20;
      6'b010101 : _zz_shift_i_3_6 = shift_i_map_21;
      6'b010110 : _zz_shift_i_3_6 = shift_i_map_22;
      6'b010111 : _zz_shift_i_3_6 = shift_i_map_23;
      6'b011000 : _zz_shift_i_3_6 = shift_i_map_24;
      6'b011001 : _zz_shift_i_3_6 = shift_i_map_25;
      6'b011010 : _zz_shift_i_3_6 = shift_i_map_26;
      6'b011011 : _zz_shift_i_3_6 = shift_i_map_27;
      6'b011100 : _zz_shift_i_3_6 = shift_i_map_28;
      6'b011101 : _zz_shift_i_3_6 = shift_i_map_29;
      6'b011110 : _zz_shift_i_3_6 = shift_i_map_30;
      6'b011111 : _zz_shift_i_3_6 = shift_i_map_31;
      6'b100000 : _zz_shift_i_3_6 = shift_i_map_32;
      6'b100001 : _zz_shift_i_3_6 = shift_i_map_33;
      6'b100010 : _zz_shift_i_3_6 = shift_i_map_34;
      6'b100011 : _zz_shift_i_3_6 = shift_i_map_35;
      6'b100100 : _zz_shift_i_3_6 = shift_i_map_36;
      6'b100101 : _zz_shift_i_3_6 = shift_i_map_37;
      6'b100110 : _zz_shift_i_3_6 = shift_i_map_38;
      6'b100111 : _zz_shift_i_3_6 = shift_i_map_39;
      6'b101000 : _zz_shift_i_3_6 = shift_i_map_40;
      6'b101001 : _zz_shift_i_3_6 = shift_i_map_41;
      6'b101010 : _zz_shift_i_3_6 = shift_i_map_42;
      6'b101011 : _zz_shift_i_3_6 = shift_i_map_43;
      6'b101100 : _zz_shift_i_3_6 = shift_i_map_44;
      6'b101101 : _zz_shift_i_3_6 = shift_i_map_45;
      6'b101110 : _zz_shift_i_3_6 = shift_i_map_46;
      6'b101111 : _zz_shift_i_3_6 = shift_i_map_47;
      6'b110000 : _zz_shift_i_3_6 = shift_i_map_48;
      6'b110001 : _zz_shift_i_3_6 = shift_i_map_49;
      6'b110010 : _zz_shift_i_3_6 = shift_i_map_50;
      6'b110011 : _zz_shift_i_3_6 = shift_i_map_51;
      6'b110100 : _zz_shift_i_3_6 = shift_i_map_52;
      6'b110101 : _zz_shift_i_3_6 = shift_i_map_53;
      6'b110110 : _zz_shift_i_3_6 = shift_i_map_54;
      6'b110111 : _zz_shift_i_3_6 = shift_i_map_55;
      6'b111000 : _zz_shift_i_3_6 = shift_i_map_56;
      6'b111001 : _zz_shift_i_3_6 = shift_i_map_57;
      6'b111010 : _zz_shift_i_3_6 = shift_i_map_58;
      6'b111011 : _zz_shift_i_3_6 = shift_i_map_59;
      6'b111100 : _zz_shift_i_3_6 = shift_i_map_60;
      6'b111101 : _zz_shift_i_3_6 = shift_i_map_61;
      6'b111110 : _zz_shift_i_3_6 = shift_i_map_62;
      default : _zz_shift_i_3_6 = shift_i_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_3_7)
      6'b000000 : _zz_shift_q_3_6 = shift_q_map_0;
      6'b000001 : _zz_shift_q_3_6 = shift_q_map_1;
      6'b000010 : _zz_shift_q_3_6 = shift_q_map_2;
      6'b000011 : _zz_shift_q_3_6 = shift_q_map_3;
      6'b000100 : _zz_shift_q_3_6 = shift_q_map_4;
      6'b000101 : _zz_shift_q_3_6 = shift_q_map_5;
      6'b000110 : _zz_shift_q_3_6 = shift_q_map_6;
      6'b000111 : _zz_shift_q_3_6 = shift_q_map_7;
      6'b001000 : _zz_shift_q_3_6 = shift_q_map_8;
      6'b001001 : _zz_shift_q_3_6 = shift_q_map_9;
      6'b001010 : _zz_shift_q_3_6 = shift_q_map_10;
      6'b001011 : _zz_shift_q_3_6 = shift_q_map_11;
      6'b001100 : _zz_shift_q_3_6 = shift_q_map_12;
      6'b001101 : _zz_shift_q_3_6 = shift_q_map_13;
      6'b001110 : _zz_shift_q_3_6 = shift_q_map_14;
      6'b001111 : _zz_shift_q_3_6 = shift_q_map_15;
      6'b010000 : _zz_shift_q_3_6 = shift_q_map_16;
      6'b010001 : _zz_shift_q_3_6 = shift_q_map_17;
      6'b010010 : _zz_shift_q_3_6 = shift_q_map_18;
      6'b010011 : _zz_shift_q_3_6 = shift_q_map_19;
      6'b010100 : _zz_shift_q_3_6 = shift_q_map_20;
      6'b010101 : _zz_shift_q_3_6 = shift_q_map_21;
      6'b010110 : _zz_shift_q_3_6 = shift_q_map_22;
      6'b010111 : _zz_shift_q_3_6 = shift_q_map_23;
      6'b011000 : _zz_shift_q_3_6 = shift_q_map_24;
      6'b011001 : _zz_shift_q_3_6 = shift_q_map_25;
      6'b011010 : _zz_shift_q_3_6 = shift_q_map_26;
      6'b011011 : _zz_shift_q_3_6 = shift_q_map_27;
      6'b011100 : _zz_shift_q_3_6 = shift_q_map_28;
      6'b011101 : _zz_shift_q_3_6 = shift_q_map_29;
      6'b011110 : _zz_shift_q_3_6 = shift_q_map_30;
      6'b011111 : _zz_shift_q_3_6 = shift_q_map_31;
      6'b100000 : _zz_shift_q_3_6 = shift_q_map_32;
      6'b100001 : _zz_shift_q_3_6 = shift_q_map_33;
      6'b100010 : _zz_shift_q_3_6 = shift_q_map_34;
      6'b100011 : _zz_shift_q_3_6 = shift_q_map_35;
      6'b100100 : _zz_shift_q_3_6 = shift_q_map_36;
      6'b100101 : _zz_shift_q_3_6 = shift_q_map_37;
      6'b100110 : _zz_shift_q_3_6 = shift_q_map_38;
      6'b100111 : _zz_shift_q_3_6 = shift_q_map_39;
      6'b101000 : _zz_shift_q_3_6 = shift_q_map_40;
      6'b101001 : _zz_shift_q_3_6 = shift_q_map_41;
      6'b101010 : _zz_shift_q_3_6 = shift_q_map_42;
      6'b101011 : _zz_shift_q_3_6 = shift_q_map_43;
      6'b101100 : _zz_shift_q_3_6 = shift_q_map_44;
      6'b101101 : _zz_shift_q_3_6 = shift_q_map_45;
      6'b101110 : _zz_shift_q_3_6 = shift_q_map_46;
      6'b101111 : _zz_shift_q_3_6 = shift_q_map_47;
      6'b110000 : _zz_shift_q_3_6 = shift_q_map_48;
      6'b110001 : _zz_shift_q_3_6 = shift_q_map_49;
      6'b110010 : _zz_shift_q_3_6 = shift_q_map_50;
      6'b110011 : _zz_shift_q_3_6 = shift_q_map_51;
      6'b110100 : _zz_shift_q_3_6 = shift_q_map_52;
      6'b110101 : _zz_shift_q_3_6 = shift_q_map_53;
      6'b110110 : _zz_shift_q_3_6 = shift_q_map_54;
      6'b110111 : _zz_shift_q_3_6 = shift_q_map_55;
      6'b111000 : _zz_shift_q_3_6 = shift_q_map_56;
      6'b111001 : _zz_shift_q_3_6 = shift_q_map_57;
      6'b111010 : _zz_shift_q_3_6 = shift_q_map_58;
      6'b111011 : _zz_shift_q_3_6 = shift_q_map_59;
      6'b111100 : _zz_shift_q_3_6 = shift_q_map_60;
      6'b111101 : _zz_shift_q_3_6 = shift_q_map_61;
      6'b111110 : _zz_shift_q_3_6 = shift_q_map_62;
      default : _zz_shift_q_3_6 = shift_q_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_4_7)
      6'b000000 : _zz_shift_i_4_6 = shift_i_map_0;
      6'b000001 : _zz_shift_i_4_6 = shift_i_map_1;
      6'b000010 : _zz_shift_i_4_6 = shift_i_map_2;
      6'b000011 : _zz_shift_i_4_6 = shift_i_map_3;
      6'b000100 : _zz_shift_i_4_6 = shift_i_map_4;
      6'b000101 : _zz_shift_i_4_6 = shift_i_map_5;
      6'b000110 : _zz_shift_i_4_6 = shift_i_map_6;
      6'b000111 : _zz_shift_i_4_6 = shift_i_map_7;
      6'b001000 : _zz_shift_i_4_6 = shift_i_map_8;
      6'b001001 : _zz_shift_i_4_6 = shift_i_map_9;
      6'b001010 : _zz_shift_i_4_6 = shift_i_map_10;
      6'b001011 : _zz_shift_i_4_6 = shift_i_map_11;
      6'b001100 : _zz_shift_i_4_6 = shift_i_map_12;
      6'b001101 : _zz_shift_i_4_6 = shift_i_map_13;
      6'b001110 : _zz_shift_i_4_6 = shift_i_map_14;
      6'b001111 : _zz_shift_i_4_6 = shift_i_map_15;
      6'b010000 : _zz_shift_i_4_6 = shift_i_map_16;
      6'b010001 : _zz_shift_i_4_6 = shift_i_map_17;
      6'b010010 : _zz_shift_i_4_6 = shift_i_map_18;
      6'b010011 : _zz_shift_i_4_6 = shift_i_map_19;
      6'b010100 : _zz_shift_i_4_6 = shift_i_map_20;
      6'b010101 : _zz_shift_i_4_6 = shift_i_map_21;
      6'b010110 : _zz_shift_i_4_6 = shift_i_map_22;
      6'b010111 : _zz_shift_i_4_6 = shift_i_map_23;
      6'b011000 : _zz_shift_i_4_6 = shift_i_map_24;
      6'b011001 : _zz_shift_i_4_6 = shift_i_map_25;
      6'b011010 : _zz_shift_i_4_6 = shift_i_map_26;
      6'b011011 : _zz_shift_i_4_6 = shift_i_map_27;
      6'b011100 : _zz_shift_i_4_6 = shift_i_map_28;
      6'b011101 : _zz_shift_i_4_6 = shift_i_map_29;
      6'b011110 : _zz_shift_i_4_6 = shift_i_map_30;
      6'b011111 : _zz_shift_i_4_6 = shift_i_map_31;
      6'b100000 : _zz_shift_i_4_6 = shift_i_map_32;
      6'b100001 : _zz_shift_i_4_6 = shift_i_map_33;
      6'b100010 : _zz_shift_i_4_6 = shift_i_map_34;
      6'b100011 : _zz_shift_i_4_6 = shift_i_map_35;
      6'b100100 : _zz_shift_i_4_6 = shift_i_map_36;
      6'b100101 : _zz_shift_i_4_6 = shift_i_map_37;
      6'b100110 : _zz_shift_i_4_6 = shift_i_map_38;
      6'b100111 : _zz_shift_i_4_6 = shift_i_map_39;
      6'b101000 : _zz_shift_i_4_6 = shift_i_map_40;
      6'b101001 : _zz_shift_i_4_6 = shift_i_map_41;
      6'b101010 : _zz_shift_i_4_6 = shift_i_map_42;
      6'b101011 : _zz_shift_i_4_6 = shift_i_map_43;
      6'b101100 : _zz_shift_i_4_6 = shift_i_map_44;
      6'b101101 : _zz_shift_i_4_6 = shift_i_map_45;
      6'b101110 : _zz_shift_i_4_6 = shift_i_map_46;
      6'b101111 : _zz_shift_i_4_6 = shift_i_map_47;
      6'b110000 : _zz_shift_i_4_6 = shift_i_map_48;
      6'b110001 : _zz_shift_i_4_6 = shift_i_map_49;
      6'b110010 : _zz_shift_i_4_6 = shift_i_map_50;
      6'b110011 : _zz_shift_i_4_6 = shift_i_map_51;
      6'b110100 : _zz_shift_i_4_6 = shift_i_map_52;
      6'b110101 : _zz_shift_i_4_6 = shift_i_map_53;
      6'b110110 : _zz_shift_i_4_6 = shift_i_map_54;
      6'b110111 : _zz_shift_i_4_6 = shift_i_map_55;
      6'b111000 : _zz_shift_i_4_6 = shift_i_map_56;
      6'b111001 : _zz_shift_i_4_6 = shift_i_map_57;
      6'b111010 : _zz_shift_i_4_6 = shift_i_map_58;
      6'b111011 : _zz_shift_i_4_6 = shift_i_map_59;
      6'b111100 : _zz_shift_i_4_6 = shift_i_map_60;
      6'b111101 : _zz_shift_i_4_6 = shift_i_map_61;
      6'b111110 : _zz_shift_i_4_6 = shift_i_map_62;
      default : _zz_shift_i_4_6 = shift_i_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_4_7)
      6'b000000 : _zz_shift_q_4_6 = shift_q_map_0;
      6'b000001 : _zz_shift_q_4_6 = shift_q_map_1;
      6'b000010 : _zz_shift_q_4_6 = shift_q_map_2;
      6'b000011 : _zz_shift_q_4_6 = shift_q_map_3;
      6'b000100 : _zz_shift_q_4_6 = shift_q_map_4;
      6'b000101 : _zz_shift_q_4_6 = shift_q_map_5;
      6'b000110 : _zz_shift_q_4_6 = shift_q_map_6;
      6'b000111 : _zz_shift_q_4_6 = shift_q_map_7;
      6'b001000 : _zz_shift_q_4_6 = shift_q_map_8;
      6'b001001 : _zz_shift_q_4_6 = shift_q_map_9;
      6'b001010 : _zz_shift_q_4_6 = shift_q_map_10;
      6'b001011 : _zz_shift_q_4_6 = shift_q_map_11;
      6'b001100 : _zz_shift_q_4_6 = shift_q_map_12;
      6'b001101 : _zz_shift_q_4_6 = shift_q_map_13;
      6'b001110 : _zz_shift_q_4_6 = shift_q_map_14;
      6'b001111 : _zz_shift_q_4_6 = shift_q_map_15;
      6'b010000 : _zz_shift_q_4_6 = shift_q_map_16;
      6'b010001 : _zz_shift_q_4_6 = shift_q_map_17;
      6'b010010 : _zz_shift_q_4_6 = shift_q_map_18;
      6'b010011 : _zz_shift_q_4_6 = shift_q_map_19;
      6'b010100 : _zz_shift_q_4_6 = shift_q_map_20;
      6'b010101 : _zz_shift_q_4_6 = shift_q_map_21;
      6'b010110 : _zz_shift_q_4_6 = shift_q_map_22;
      6'b010111 : _zz_shift_q_4_6 = shift_q_map_23;
      6'b011000 : _zz_shift_q_4_6 = shift_q_map_24;
      6'b011001 : _zz_shift_q_4_6 = shift_q_map_25;
      6'b011010 : _zz_shift_q_4_6 = shift_q_map_26;
      6'b011011 : _zz_shift_q_4_6 = shift_q_map_27;
      6'b011100 : _zz_shift_q_4_6 = shift_q_map_28;
      6'b011101 : _zz_shift_q_4_6 = shift_q_map_29;
      6'b011110 : _zz_shift_q_4_6 = shift_q_map_30;
      6'b011111 : _zz_shift_q_4_6 = shift_q_map_31;
      6'b100000 : _zz_shift_q_4_6 = shift_q_map_32;
      6'b100001 : _zz_shift_q_4_6 = shift_q_map_33;
      6'b100010 : _zz_shift_q_4_6 = shift_q_map_34;
      6'b100011 : _zz_shift_q_4_6 = shift_q_map_35;
      6'b100100 : _zz_shift_q_4_6 = shift_q_map_36;
      6'b100101 : _zz_shift_q_4_6 = shift_q_map_37;
      6'b100110 : _zz_shift_q_4_6 = shift_q_map_38;
      6'b100111 : _zz_shift_q_4_6 = shift_q_map_39;
      6'b101000 : _zz_shift_q_4_6 = shift_q_map_40;
      6'b101001 : _zz_shift_q_4_6 = shift_q_map_41;
      6'b101010 : _zz_shift_q_4_6 = shift_q_map_42;
      6'b101011 : _zz_shift_q_4_6 = shift_q_map_43;
      6'b101100 : _zz_shift_q_4_6 = shift_q_map_44;
      6'b101101 : _zz_shift_q_4_6 = shift_q_map_45;
      6'b101110 : _zz_shift_q_4_6 = shift_q_map_46;
      6'b101111 : _zz_shift_q_4_6 = shift_q_map_47;
      6'b110000 : _zz_shift_q_4_6 = shift_q_map_48;
      6'b110001 : _zz_shift_q_4_6 = shift_q_map_49;
      6'b110010 : _zz_shift_q_4_6 = shift_q_map_50;
      6'b110011 : _zz_shift_q_4_6 = shift_q_map_51;
      6'b110100 : _zz_shift_q_4_6 = shift_q_map_52;
      6'b110101 : _zz_shift_q_4_6 = shift_q_map_53;
      6'b110110 : _zz_shift_q_4_6 = shift_q_map_54;
      6'b110111 : _zz_shift_q_4_6 = shift_q_map_55;
      6'b111000 : _zz_shift_q_4_6 = shift_q_map_56;
      6'b111001 : _zz_shift_q_4_6 = shift_q_map_57;
      6'b111010 : _zz_shift_q_4_6 = shift_q_map_58;
      6'b111011 : _zz_shift_q_4_6 = shift_q_map_59;
      6'b111100 : _zz_shift_q_4_6 = shift_q_map_60;
      6'b111101 : _zz_shift_q_4_6 = shift_q_map_61;
      6'b111110 : _zz_shift_q_4_6 = shift_q_map_62;
      default : _zz_shift_q_4_6 = shift_q_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_5_7)
      6'b000000 : _zz_shift_i_5_6 = shift_i_map_0;
      6'b000001 : _zz_shift_i_5_6 = shift_i_map_1;
      6'b000010 : _zz_shift_i_5_6 = shift_i_map_2;
      6'b000011 : _zz_shift_i_5_6 = shift_i_map_3;
      6'b000100 : _zz_shift_i_5_6 = shift_i_map_4;
      6'b000101 : _zz_shift_i_5_6 = shift_i_map_5;
      6'b000110 : _zz_shift_i_5_6 = shift_i_map_6;
      6'b000111 : _zz_shift_i_5_6 = shift_i_map_7;
      6'b001000 : _zz_shift_i_5_6 = shift_i_map_8;
      6'b001001 : _zz_shift_i_5_6 = shift_i_map_9;
      6'b001010 : _zz_shift_i_5_6 = shift_i_map_10;
      6'b001011 : _zz_shift_i_5_6 = shift_i_map_11;
      6'b001100 : _zz_shift_i_5_6 = shift_i_map_12;
      6'b001101 : _zz_shift_i_5_6 = shift_i_map_13;
      6'b001110 : _zz_shift_i_5_6 = shift_i_map_14;
      6'b001111 : _zz_shift_i_5_6 = shift_i_map_15;
      6'b010000 : _zz_shift_i_5_6 = shift_i_map_16;
      6'b010001 : _zz_shift_i_5_6 = shift_i_map_17;
      6'b010010 : _zz_shift_i_5_6 = shift_i_map_18;
      6'b010011 : _zz_shift_i_5_6 = shift_i_map_19;
      6'b010100 : _zz_shift_i_5_6 = shift_i_map_20;
      6'b010101 : _zz_shift_i_5_6 = shift_i_map_21;
      6'b010110 : _zz_shift_i_5_6 = shift_i_map_22;
      6'b010111 : _zz_shift_i_5_6 = shift_i_map_23;
      6'b011000 : _zz_shift_i_5_6 = shift_i_map_24;
      6'b011001 : _zz_shift_i_5_6 = shift_i_map_25;
      6'b011010 : _zz_shift_i_5_6 = shift_i_map_26;
      6'b011011 : _zz_shift_i_5_6 = shift_i_map_27;
      6'b011100 : _zz_shift_i_5_6 = shift_i_map_28;
      6'b011101 : _zz_shift_i_5_6 = shift_i_map_29;
      6'b011110 : _zz_shift_i_5_6 = shift_i_map_30;
      6'b011111 : _zz_shift_i_5_6 = shift_i_map_31;
      6'b100000 : _zz_shift_i_5_6 = shift_i_map_32;
      6'b100001 : _zz_shift_i_5_6 = shift_i_map_33;
      6'b100010 : _zz_shift_i_5_6 = shift_i_map_34;
      6'b100011 : _zz_shift_i_5_6 = shift_i_map_35;
      6'b100100 : _zz_shift_i_5_6 = shift_i_map_36;
      6'b100101 : _zz_shift_i_5_6 = shift_i_map_37;
      6'b100110 : _zz_shift_i_5_6 = shift_i_map_38;
      6'b100111 : _zz_shift_i_5_6 = shift_i_map_39;
      6'b101000 : _zz_shift_i_5_6 = shift_i_map_40;
      6'b101001 : _zz_shift_i_5_6 = shift_i_map_41;
      6'b101010 : _zz_shift_i_5_6 = shift_i_map_42;
      6'b101011 : _zz_shift_i_5_6 = shift_i_map_43;
      6'b101100 : _zz_shift_i_5_6 = shift_i_map_44;
      6'b101101 : _zz_shift_i_5_6 = shift_i_map_45;
      6'b101110 : _zz_shift_i_5_6 = shift_i_map_46;
      6'b101111 : _zz_shift_i_5_6 = shift_i_map_47;
      6'b110000 : _zz_shift_i_5_6 = shift_i_map_48;
      6'b110001 : _zz_shift_i_5_6 = shift_i_map_49;
      6'b110010 : _zz_shift_i_5_6 = shift_i_map_50;
      6'b110011 : _zz_shift_i_5_6 = shift_i_map_51;
      6'b110100 : _zz_shift_i_5_6 = shift_i_map_52;
      6'b110101 : _zz_shift_i_5_6 = shift_i_map_53;
      6'b110110 : _zz_shift_i_5_6 = shift_i_map_54;
      6'b110111 : _zz_shift_i_5_6 = shift_i_map_55;
      6'b111000 : _zz_shift_i_5_6 = shift_i_map_56;
      6'b111001 : _zz_shift_i_5_6 = shift_i_map_57;
      6'b111010 : _zz_shift_i_5_6 = shift_i_map_58;
      6'b111011 : _zz_shift_i_5_6 = shift_i_map_59;
      6'b111100 : _zz_shift_i_5_6 = shift_i_map_60;
      6'b111101 : _zz_shift_i_5_6 = shift_i_map_61;
      6'b111110 : _zz_shift_i_5_6 = shift_i_map_62;
      default : _zz_shift_i_5_6 = shift_i_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_5_7)
      6'b000000 : _zz_shift_q_5_6 = shift_q_map_0;
      6'b000001 : _zz_shift_q_5_6 = shift_q_map_1;
      6'b000010 : _zz_shift_q_5_6 = shift_q_map_2;
      6'b000011 : _zz_shift_q_5_6 = shift_q_map_3;
      6'b000100 : _zz_shift_q_5_6 = shift_q_map_4;
      6'b000101 : _zz_shift_q_5_6 = shift_q_map_5;
      6'b000110 : _zz_shift_q_5_6 = shift_q_map_6;
      6'b000111 : _zz_shift_q_5_6 = shift_q_map_7;
      6'b001000 : _zz_shift_q_5_6 = shift_q_map_8;
      6'b001001 : _zz_shift_q_5_6 = shift_q_map_9;
      6'b001010 : _zz_shift_q_5_6 = shift_q_map_10;
      6'b001011 : _zz_shift_q_5_6 = shift_q_map_11;
      6'b001100 : _zz_shift_q_5_6 = shift_q_map_12;
      6'b001101 : _zz_shift_q_5_6 = shift_q_map_13;
      6'b001110 : _zz_shift_q_5_6 = shift_q_map_14;
      6'b001111 : _zz_shift_q_5_6 = shift_q_map_15;
      6'b010000 : _zz_shift_q_5_6 = shift_q_map_16;
      6'b010001 : _zz_shift_q_5_6 = shift_q_map_17;
      6'b010010 : _zz_shift_q_5_6 = shift_q_map_18;
      6'b010011 : _zz_shift_q_5_6 = shift_q_map_19;
      6'b010100 : _zz_shift_q_5_6 = shift_q_map_20;
      6'b010101 : _zz_shift_q_5_6 = shift_q_map_21;
      6'b010110 : _zz_shift_q_5_6 = shift_q_map_22;
      6'b010111 : _zz_shift_q_5_6 = shift_q_map_23;
      6'b011000 : _zz_shift_q_5_6 = shift_q_map_24;
      6'b011001 : _zz_shift_q_5_6 = shift_q_map_25;
      6'b011010 : _zz_shift_q_5_6 = shift_q_map_26;
      6'b011011 : _zz_shift_q_5_6 = shift_q_map_27;
      6'b011100 : _zz_shift_q_5_6 = shift_q_map_28;
      6'b011101 : _zz_shift_q_5_6 = shift_q_map_29;
      6'b011110 : _zz_shift_q_5_6 = shift_q_map_30;
      6'b011111 : _zz_shift_q_5_6 = shift_q_map_31;
      6'b100000 : _zz_shift_q_5_6 = shift_q_map_32;
      6'b100001 : _zz_shift_q_5_6 = shift_q_map_33;
      6'b100010 : _zz_shift_q_5_6 = shift_q_map_34;
      6'b100011 : _zz_shift_q_5_6 = shift_q_map_35;
      6'b100100 : _zz_shift_q_5_6 = shift_q_map_36;
      6'b100101 : _zz_shift_q_5_6 = shift_q_map_37;
      6'b100110 : _zz_shift_q_5_6 = shift_q_map_38;
      6'b100111 : _zz_shift_q_5_6 = shift_q_map_39;
      6'b101000 : _zz_shift_q_5_6 = shift_q_map_40;
      6'b101001 : _zz_shift_q_5_6 = shift_q_map_41;
      6'b101010 : _zz_shift_q_5_6 = shift_q_map_42;
      6'b101011 : _zz_shift_q_5_6 = shift_q_map_43;
      6'b101100 : _zz_shift_q_5_6 = shift_q_map_44;
      6'b101101 : _zz_shift_q_5_6 = shift_q_map_45;
      6'b101110 : _zz_shift_q_5_6 = shift_q_map_46;
      6'b101111 : _zz_shift_q_5_6 = shift_q_map_47;
      6'b110000 : _zz_shift_q_5_6 = shift_q_map_48;
      6'b110001 : _zz_shift_q_5_6 = shift_q_map_49;
      6'b110010 : _zz_shift_q_5_6 = shift_q_map_50;
      6'b110011 : _zz_shift_q_5_6 = shift_q_map_51;
      6'b110100 : _zz_shift_q_5_6 = shift_q_map_52;
      6'b110101 : _zz_shift_q_5_6 = shift_q_map_53;
      6'b110110 : _zz_shift_q_5_6 = shift_q_map_54;
      6'b110111 : _zz_shift_q_5_6 = shift_q_map_55;
      6'b111000 : _zz_shift_q_5_6 = shift_q_map_56;
      6'b111001 : _zz_shift_q_5_6 = shift_q_map_57;
      6'b111010 : _zz_shift_q_5_6 = shift_q_map_58;
      6'b111011 : _zz_shift_q_5_6 = shift_q_map_59;
      6'b111100 : _zz_shift_q_5_6 = shift_q_map_60;
      6'b111101 : _zz_shift_q_5_6 = shift_q_map_61;
      6'b111110 : _zz_shift_q_5_6 = shift_q_map_62;
      default : _zz_shift_q_5_6 = shift_q_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_6_7)
      6'b000000 : _zz_shift_i_6_6 = shift_i_map_0;
      6'b000001 : _zz_shift_i_6_6 = shift_i_map_1;
      6'b000010 : _zz_shift_i_6_6 = shift_i_map_2;
      6'b000011 : _zz_shift_i_6_6 = shift_i_map_3;
      6'b000100 : _zz_shift_i_6_6 = shift_i_map_4;
      6'b000101 : _zz_shift_i_6_6 = shift_i_map_5;
      6'b000110 : _zz_shift_i_6_6 = shift_i_map_6;
      6'b000111 : _zz_shift_i_6_6 = shift_i_map_7;
      6'b001000 : _zz_shift_i_6_6 = shift_i_map_8;
      6'b001001 : _zz_shift_i_6_6 = shift_i_map_9;
      6'b001010 : _zz_shift_i_6_6 = shift_i_map_10;
      6'b001011 : _zz_shift_i_6_6 = shift_i_map_11;
      6'b001100 : _zz_shift_i_6_6 = shift_i_map_12;
      6'b001101 : _zz_shift_i_6_6 = shift_i_map_13;
      6'b001110 : _zz_shift_i_6_6 = shift_i_map_14;
      6'b001111 : _zz_shift_i_6_6 = shift_i_map_15;
      6'b010000 : _zz_shift_i_6_6 = shift_i_map_16;
      6'b010001 : _zz_shift_i_6_6 = shift_i_map_17;
      6'b010010 : _zz_shift_i_6_6 = shift_i_map_18;
      6'b010011 : _zz_shift_i_6_6 = shift_i_map_19;
      6'b010100 : _zz_shift_i_6_6 = shift_i_map_20;
      6'b010101 : _zz_shift_i_6_6 = shift_i_map_21;
      6'b010110 : _zz_shift_i_6_6 = shift_i_map_22;
      6'b010111 : _zz_shift_i_6_6 = shift_i_map_23;
      6'b011000 : _zz_shift_i_6_6 = shift_i_map_24;
      6'b011001 : _zz_shift_i_6_6 = shift_i_map_25;
      6'b011010 : _zz_shift_i_6_6 = shift_i_map_26;
      6'b011011 : _zz_shift_i_6_6 = shift_i_map_27;
      6'b011100 : _zz_shift_i_6_6 = shift_i_map_28;
      6'b011101 : _zz_shift_i_6_6 = shift_i_map_29;
      6'b011110 : _zz_shift_i_6_6 = shift_i_map_30;
      6'b011111 : _zz_shift_i_6_6 = shift_i_map_31;
      6'b100000 : _zz_shift_i_6_6 = shift_i_map_32;
      6'b100001 : _zz_shift_i_6_6 = shift_i_map_33;
      6'b100010 : _zz_shift_i_6_6 = shift_i_map_34;
      6'b100011 : _zz_shift_i_6_6 = shift_i_map_35;
      6'b100100 : _zz_shift_i_6_6 = shift_i_map_36;
      6'b100101 : _zz_shift_i_6_6 = shift_i_map_37;
      6'b100110 : _zz_shift_i_6_6 = shift_i_map_38;
      6'b100111 : _zz_shift_i_6_6 = shift_i_map_39;
      6'b101000 : _zz_shift_i_6_6 = shift_i_map_40;
      6'b101001 : _zz_shift_i_6_6 = shift_i_map_41;
      6'b101010 : _zz_shift_i_6_6 = shift_i_map_42;
      6'b101011 : _zz_shift_i_6_6 = shift_i_map_43;
      6'b101100 : _zz_shift_i_6_6 = shift_i_map_44;
      6'b101101 : _zz_shift_i_6_6 = shift_i_map_45;
      6'b101110 : _zz_shift_i_6_6 = shift_i_map_46;
      6'b101111 : _zz_shift_i_6_6 = shift_i_map_47;
      6'b110000 : _zz_shift_i_6_6 = shift_i_map_48;
      6'b110001 : _zz_shift_i_6_6 = shift_i_map_49;
      6'b110010 : _zz_shift_i_6_6 = shift_i_map_50;
      6'b110011 : _zz_shift_i_6_6 = shift_i_map_51;
      6'b110100 : _zz_shift_i_6_6 = shift_i_map_52;
      6'b110101 : _zz_shift_i_6_6 = shift_i_map_53;
      6'b110110 : _zz_shift_i_6_6 = shift_i_map_54;
      6'b110111 : _zz_shift_i_6_6 = shift_i_map_55;
      6'b111000 : _zz_shift_i_6_6 = shift_i_map_56;
      6'b111001 : _zz_shift_i_6_6 = shift_i_map_57;
      6'b111010 : _zz_shift_i_6_6 = shift_i_map_58;
      6'b111011 : _zz_shift_i_6_6 = shift_i_map_59;
      6'b111100 : _zz_shift_i_6_6 = shift_i_map_60;
      6'b111101 : _zz_shift_i_6_6 = shift_i_map_61;
      6'b111110 : _zz_shift_i_6_6 = shift_i_map_62;
      default : _zz_shift_i_6_6 = shift_i_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_6_7)
      6'b000000 : _zz_shift_q_6_6 = shift_q_map_0;
      6'b000001 : _zz_shift_q_6_6 = shift_q_map_1;
      6'b000010 : _zz_shift_q_6_6 = shift_q_map_2;
      6'b000011 : _zz_shift_q_6_6 = shift_q_map_3;
      6'b000100 : _zz_shift_q_6_6 = shift_q_map_4;
      6'b000101 : _zz_shift_q_6_6 = shift_q_map_5;
      6'b000110 : _zz_shift_q_6_6 = shift_q_map_6;
      6'b000111 : _zz_shift_q_6_6 = shift_q_map_7;
      6'b001000 : _zz_shift_q_6_6 = shift_q_map_8;
      6'b001001 : _zz_shift_q_6_6 = shift_q_map_9;
      6'b001010 : _zz_shift_q_6_6 = shift_q_map_10;
      6'b001011 : _zz_shift_q_6_6 = shift_q_map_11;
      6'b001100 : _zz_shift_q_6_6 = shift_q_map_12;
      6'b001101 : _zz_shift_q_6_6 = shift_q_map_13;
      6'b001110 : _zz_shift_q_6_6 = shift_q_map_14;
      6'b001111 : _zz_shift_q_6_6 = shift_q_map_15;
      6'b010000 : _zz_shift_q_6_6 = shift_q_map_16;
      6'b010001 : _zz_shift_q_6_6 = shift_q_map_17;
      6'b010010 : _zz_shift_q_6_6 = shift_q_map_18;
      6'b010011 : _zz_shift_q_6_6 = shift_q_map_19;
      6'b010100 : _zz_shift_q_6_6 = shift_q_map_20;
      6'b010101 : _zz_shift_q_6_6 = shift_q_map_21;
      6'b010110 : _zz_shift_q_6_6 = shift_q_map_22;
      6'b010111 : _zz_shift_q_6_6 = shift_q_map_23;
      6'b011000 : _zz_shift_q_6_6 = shift_q_map_24;
      6'b011001 : _zz_shift_q_6_6 = shift_q_map_25;
      6'b011010 : _zz_shift_q_6_6 = shift_q_map_26;
      6'b011011 : _zz_shift_q_6_6 = shift_q_map_27;
      6'b011100 : _zz_shift_q_6_6 = shift_q_map_28;
      6'b011101 : _zz_shift_q_6_6 = shift_q_map_29;
      6'b011110 : _zz_shift_q_6_6 = shift_q_map_30;
      6'b011111 : _zz_shift_q_6_6 = shift_q_map_31;
      6'b100000 : _zz_shift_q_6_6 = shift_q_map_32;
      6'b100001 : _zz_shift_q_6_6 = shift_q_map_33;
      6'b100010 : _zz_shift_q_6_6 = shift_q_map_34;
      6'b100011 : _zz_shift_q_6_6 = shift_q_map_35;
      6'b100100 : _zz_shift_q_6_6 = shift_q_map_36;
      6'b100101 : _zz_shift_q_6_6 = shift_q_map_37;
      6'b100110 : _zz_shift_q_6_6 = shift_q_map_38;
      6'b100111 : _zz_shift_q_6_6 = shift_q_map_39;
      6'b101000 : _zz_shift_q_6_6 = shift_q_map_40;
      6'b101001 : _zz_shift_q_6_6 = shift_q_map_41;
      6'b101010 : _zz_shift_q_6_6 = shift_q_map_42;
      6'b101011 : _zz_shift_q_6_6 = shift_q_map_43;
      6'b101100 : _zz_shift_q_6_6 = shift_q_map_44;
      6'b101101 : _zz_shift_q_6_6 = shift_q_map_45;
      6'b101110 : _zz_shift_q_6_6 = shift_q_map_46;
      6'b101111 : _zz_shift_q_6_6 = shift_q_map_47;
      6'b110000 : _zz_shift_q_6_6 = shift_q_map_48;
      6'b110001 : _zz_shift_q_6_6 = shift_q_map_49;
      6'b110010 : _zz_shift_q_6_6 = shift_q_map_50;
      6'b110011 : _zz_shift_q_6_6 = shift_q_map_51;
      6'b110100 : _zz_shift_q_6_6 = shift_q_map_52;
      6'b110101 : _zz_shift_q_6_6 = shift_q_map_53;
      6'b110110 : _zz_shift_q_6_6 = shift_q_map_54;
      6'b110111 : _zz_shift_q_6_6 = shift_q_map_55;
      6'b111000 : _zz_shift_q_6_6 = shift_q_map_56;
      6'b111001 : _zz_shift_q_6_6 = shift_q_map_57;
      6'b111010 : _zz_shift_q_6_6 = shift_q_map_58;
      6'b111011 : _zz_shift_q_6_6 = shift_q_map_59;
      6'b111100 : _zz_shift_q_6_6 = shift_q_map_60;
      6'b111101 : _zz_shift_q_6_6 = shift_q_map_61;
      6'b111110 : _zz_shift_q_6_6 = shift_q_map_62;
      default : _zz_shift_q_6_6 = shift_q_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_7_7)
      6'b000000 : _zz_shift_i_7_6 = shift_i_map_0;
      6'b000001 : _zz_shift_i_7_6 = shift_i_map_1;
      6'b000010 : _zz_shift_i_7_6 = shift_i_map_2;
      6'b000011 : _zz_shift_i_7_6 = shift_i_map_3;
      6'b000100 : _zz_shift_i_7_6 = shift_i_map_4;
      6'b000101 : _zz_shift_i_7_6 = shift_i_map_5;
      6'b000110 : _zz_shift_i_7_6 = shift_i_map_6;
      6'b000111 : _zz_shift_i_7_6 = shift_i_map_7;
      6'b001000 : _zz_shift_i_7_6 = shift_i_map_8;
      6'b001001 : _zz_shift_i_7_6 = shift_i_map_9;
      6'b001010 : _zz_shift_i_7_6 = shift_i_map_10;
      6'b001011 : _zz_shift_i_7_6 = shift_i_map_11;
      6'b001100 : _zz_shift_i_7_6 = shift_i_map_12;
      6'b001101 : _zz_shift_i_7_6 = shift_i_map_13;
      6'b001110 : _zz_shift_i_7_6 = shift_i_map_14;
      6'b001111 : _zz_shift_i_7_6 = shift_i_map_15;
      6'b010000 : _zz_shift_i_7_6 = shift_i_map_16;
      6'b010001 : _zz_shift_i_7_6 = shift_i_map_17;
      6'b010010 : _zz_shift_i_7_6 = shift_i_map_18;
      6'b010011 : _zz_shift_i_7_6 = shift_i_map_19;
      6'b010100 : _zz_shift_i_7_6 = shift_i_map_20;
      6'b010101 : _zz_shift_i_7_6 = shift_i_map_21;
      6'b010110 : _zz_shift_i_7_6 = shift_i_map_22;
      6'b010111 : _zz_shift_i_7_6 = shift_i_map_23;
      6'b011000 : _zz_shift_i_7_6 = shift_i_map_24;
      6'b011001 : _zz_shift_i_7_6 = shift_i_map_25;
      6'b011010 : _zz_shift_i_7_6 = shift_i_map_26;
      6'b011011 : _zz_shift_i_7_6 = shift_i_map_27;
      6'b011100 : _zz_shift_i_7_6 = shift_i_map_28;
      6'b011101 : _zz_shift_i_7_6 = shift_i_map_29;
      6'b011110 : _zz_shift_i_7_6 = shift_i_map_30;
      6'b011111 : _zz_shift_i_7_6 = shift_i_map_31;
      6'b100000 : _zz_shift_i_7_6 = shift_i_map_32;
      6'b100001 : _zz_shift_i_7_6 = shift_i_map_33;
      6'b100010 : _zz_shift_i_7_6 = shift_i_map_34;
      6'b100011 : _zz_shift_i_7_6 = shift_i_map_35;
      6'b100100 : _zz_shift_i_7_6 = shift_i_map_36;
      6'b100101 : _zz_shift_i_7_6 = shift_i_map_37;
      6'b100110 : _zz_shift_i_7_6 = shift_i_map_38;
      6'b100111 : _zz_shift_i_7_6 = shift_i_map_39;
      6'b101000 : _zz_shift_i_7_6 = shift_i_map_40;
      6'b101001 : _zz_shift_i_7_6 = shift_i_map_41;
      6'b101010 : _zz_shift_i_7_6 = shift_i_map_42;
      6'b101011 : _zz_shift_i_7_6 = shift_i_map_43;
      6'b101100 : _zz_shift_i_7_6 = shift_i_map_44;
      6'b101101 : _zz_shift_i_7_6 = shift_i_map_45;
      6'b101110 : _zz_shift_i_7_6 = shift_i_map_46;
      6'b101111 : _zz_shift_i_7_6 = shift_i_map_47;
      6'b110000 : _zz_shift_i_7_6 = shift_i_map_48;
      6'b110001 : _zz_shift_i_7_6 = shift_i_map_49;
      6'b110010 : _zz_shift_i_7_6 = shift_i_map_50;
      6'b110011 : _zz_shift_i_7_6 = shift_i_map_51;
      6'b110100 : _zz_shift_i_7_6 = shift_i_map_52;
      6'b110101 : _zz_shift_i_7_6 = shift_i_map_53;
      6'b110110 : _zz_shift_i_7_6 = shift_i_map_54;
      6'b110111 : _zz_shift_i_7_6 = shift_i_map_55;
      6'b111000 : _zz_shift_i_7_6 = shift_i_map_56;
      6'b111001 : _zz_shift_i_7_6 = shift_i_map_57;
      6'b111010 : _zz_shift_i_7_6 = shift_i_map_58;
      6'b111011 : _zz_shift_i_7_6 = shift_i_map_59;
      6'b111100 : _zz_shift_i_7_6 = shift_i_map_60;
      6'b111101 : _zz_shift_i_7_6 = shift_i_map_61;
      6'b111110 : _zz_shift_i_7_6 = shift_i_map_62;
      default : _zz_shift_i_7_6 = shift_i_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_7_7)
      6'b000000 : _zz_shift_q_7_6 = shift_q_map_0;
      6'b000001 : _zz_shift_q_7_6 = shift_q_map_1;
      6'b000010 : _zz_shift_q_7_6 = shift_q_map_2;
      6'b000011 : _zz_shift_q_7_6 = shift_q_map_3;
      6'b000100 : _zz_shift_q_7_6 = shift_q_map_4;
      6'b000101 : _zz_shift_q_7_6 = shift_q_map_5;
      6'b000110 : _zz_shift_q_7_6 = shift_q_map_6;
      6'b000111 : _zz_shift_q_7_6 = shift_q_map_7;
      6'b001000 : _zz_shift_q_7_6 = shift_q_map_8;
      6'b001001 : _zz_shift_q_7_6 = shift_q_map_9;
      6'b001010 : _zz_shift_q_7_6 = shift_q_map_10;
      6'b001011 : _zz_shift_q_7_6 = shift_q_map_11;
      6'b001100 : _zz_shift_q_7_6 = shift_q_map_12;
      6'b001101 : _zz_shift_q_7_6 = shift_q_map_13;
      6'b001110 : _zz_shift_q_7_6 = shift_q_map_14;
      6'b001111 : _zz_shift_q_7_6 = shift_q_map_15;
      6'b010000 : _zz_shift_q_7_6 = shift_q_map_16;
      6'b010001 : _zz_shift_q_7_6 = shift_q_map_17;
      6'b010010 : _zz_shift_q_7_6 = shift_q_map_18;
      6'b010011 : _zz_shift_q_7_6 = shift_q_map_19;
      6'b010100 : _zz_shift_q_7_6 = shift_q_map_20;
      6'b010101 : _zz_shift_q_7_6 = shift_q_map_21;
      6'b010110 : _zz_shift_q_7_6 = shift_q_map_22;
      6'b010111 : _zz_shift_q_7_6 = shift_q_map_23;
      6'b011000 : _zz_shift_q_7_6 = shift_q_map_24;
      6'b011001 : _zz_shift_q_7_6 = shift_q_map_25;
      6'b011010 : _zz_shift_q_7_6 = shift_q_map_26;
      6'b011011 : _zz_shift_q_7_6 = shift_q_map_27;
      6'b011100 : _zz_shift_q_7_6 = shift_q_map_28;
      6'b011101 : _zz_shift_q_7_6 = shift_q_map_29;
      6'b011110 : _zz_shift_q_7_6 = shift_q_map_30;
      6'b011111 : _zz_shift_q_7_6 = shift_q_map_31;
      6'b100000 : _zz_shift_q_7_6 = shift_q_map_32;
      6'b100001 : _zz_shift_q_7_6 = shift_q_map_33;
      6'b100010 : _zz_shift_q_7_6 = shift_q_map_34;
      6'b100011 : _zz_shift_q_7_6 = shift_q_map_35;
      6'b100100 : _zz_shift_q_7_6 = shift_q_map_36;
      6'b100101 : _zz_shift_q_7_6 = shift_q_map_37;
      6'b100110 : _zz_shift_q_7_6 = shift_q_map_38;
      6'b100111 : _zz_shift_q_7_6 = shift_q_map_39;
      6'b101000 : _zz_shift_q_7_6 = shift_q_map_40;
      6'b101001 : _zz_shift_q_7_6 = shift_q_map_41;
      6'b101010 : _zz_shift_q_7_6 = shift_q_map_42;
      6'b101011 : _zz_shift_q_7_6 = shift_q_map_43;
      6'b101100 : _zz_shift_q_7_6 = shift_q_map_44;
      6'b101101 : _zz_shift_q_7_6 = shift_q_map_45;
      6'b101110 : _zz_shift_q_7_6 = shift_q_map_46;
      6'b101111 : _zz_shift_q_7_6 = shift_q_map_47;
      6'b110000 : _zz_shift_q_7_6 = shift_q_map_48;
      6'b110001 : _zz_shift_q_7_6 = shift_q_map_49;
      6'b110010 : _zz_shift_q_7_6 = shift_q_map_50;
      6'b110011 : _zz_shift_q_7_6 = shift_q_map_51;
      6'b110100 : _zz_shift_q_7_6 = shift_q_map_52;
      6'b110101 : _zz_shift_q_7_6 = shift_q_map_53;
      6'b110110 : _zz_shift_q_7_6 = shift_q_map_54;
      6'b110111 : _zz_shift_q_7_6 = shift_q_map_55;
      6'b111000 : _zz_shift_q_7_6 = shift_q_map_56;
      6'b111001 : _zz_shift_q_7_6 = shift_q_map_57;
      6'b111010 : _zz_shift_q_7_6 = shift_q_map_58;
      6'b111011 : _zz_shift_q_7_6 = shift_q_map_59;
      6'b111100 : _zz_shift_q_7_6 = shift_q_map_60;
      6'b111101 : _zz_shift_q_7_6 = shift_q_map_61;
      6'b111110 : _zz_shift_q_7_6 = shift_q_map_62;
      default : _zz_shift_q_7_6 = shift_q_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_0_9)
      6'b000000 : _zz_shift_i_0_8 = shift_i_map_0;
      6'b000001 : _zz_shift_i_0_8 = shift_i_map_1;
      6'b000010 : _zz_shift_i_0_8 = shift_i_map_2;
      6'b000011 : _zz_shift_i_0_8 = shift_i_map_3;
      6'b000100 : _zz_shift_i_0_8 = shift_i_map_4;
      6'b000101 : _zz_shift_i_0_8 = shift_i_map_5;
      6'b000110 : _zz_shift_i_0_8 = shift_i_map_6;
      6'b000111 : _zz_shift_i_0_8 = shift_i_map_7;
      6'b001000 : _zz_shift_i_0_8 = shift_i_map_8;
      6'b001001 : _zz_shift_i_0_8 = shift_i_map_9;
      6'b001010 : _zz_shift_i_0_8 = shift_i_map_10;
      6'b001011 : _zz_shift_i_0_8 = shift_i_map_11;
      6'b001100 : _zz_shift_i_0_8 = shift_i_map_12;
      6'b001101 : _zz_shift_i_0_8 = shift_i_map_13;
      6'b001110 : _zz_shift_i_0_8 = shift_i_map_14;
      6'b001111 : _zz_shift_i_0_8 = shift_i_map_15;
      6'b010000 : _zz_shift_i_0_8 = shift_i_map_16;
      6'b010001 : _zz_shift_i_0_8 = shift_i_map_17;
      6'b010010 : _zz_shift_i_0_8 = shift_i_map_18;
      6'b010011 : _zz_shift_i_0_8 = shift_i_map_19;
      6'b010100 : _zz_shift_i_0_8 = shift_i_map_20;
      6'b010101 : _zz_shift_i_0_8 = shift_i_map_21;
      6'b010110 : _zz_shift_i_0_8 = shift_i_map_22;
      6'b010111 : _zz_shift_i_0_8 = shift_i_map_23;
      6'b011000 : _zz_shift_i_0_8 = shift_i_map_24;
      6'b011001 : _zz_shift_i_0_8 = shift_i_map_25;
      6'b011010 : _zz_shift_i_0_8 = shift_i_map_26;
      6'b011011 : _zz_shift_i_0_8 = shift_i_map_27;
      6'b011100 : _zz_shift_i_0_8 = shift_i_map_28;
      6'b011101 : _zz_shift_i_0_8 = shift_i_map_29;
      6'b011110 : _zz_shift_i_0_8 = shift_i_map_30;
      6'b011111 : _zz_shift_i_0_8 = shift_i_map_31;
      6'b100000 : _zz_shift_i_0_8 = shift_i_map_32;
      6'b100001 : _zz_shift_i_0_8 = shift_i_map_33;
      6'b100010 : _zz_shift_i_0_8 = shift_i_map_34;
      6'b100011 : _zz_shift_i_0_8 = shift_i_map_35;
      6'b100100 : _zz_shift_i_0_8 = shift_i_map_36;
      6'b100101 : _zz_shift_i_0_8 = shift_i_map_37;
      6'b100110 : _zz_shift_i_0_8 = shift_i_map_38;
      6'b100111 : _zz_shift_i_0_8 = shift_i_map_39;
      6'b101000 : _zz_shift_i_0_8 = shift_i_map_40;
      6'b101001 : _zz_shift_i_0_8 = shift_i_map_41;
      6'b101010 : _zz_shift_i_0_8 = shift_i_map_42;
      6'b101011 : _zz_shift_i_0_8 = shift_i_map_43;
      6'b101100 : _zz_shift_i_0_8 = shift_i_map_44;
      6'b101101 : _zz_shift_i_0_8 = shift_i_map_45;
      6'b101110 : _zz_shift_i_0_8 = shift_i_map_46;
      6'b101111 : _zz_shift_i_0_8 = shift_i_map_47;
      6'b110000 : _zz_shift_i_0_8 = shift_i_map_48;
      6'b110001 : _zz_shift_i_0_8 = shift_i_map_49;
      6'b110010 : _zz_shift_i_0_8 = shift_i_map_50;
      6'b110011 : _zz_shift_i_0_8 = shift_i_map_51;
      6'b110100 : _zz_shift_i_0_8 = shift_i_map_52;
      6'b110101 : _zz_shift_i_0_8 = shift_i_map_53;
      6'b110110 : _zz_shift_i_0_8 = shift_i_map_54;
      6'b110111 : _zz_shift_i_0_8 = shift_i_map_55;
      6'b111000 : _zz_shift_i_0_8 = shift_i_map_56;
      6'b111001 : _zz_shift_i_0_8 = shift_i_map_57;
      6'b111010 : _zz_shift_i_0_8 = shift_i_map_58;
      6'b111011 : _zz_shift_i_0_8 = shift_i_map_59;
      6'b111100 : _zz_shift_i_0_8 = shift_i_map_60;
      6'b111101 : _zz_shift_i_0_8 = shift_i_map_61;
      6'b111110 : _zz_shift_i_0_8 = shift_i_map_62;
      default : _zz_shift_i_0_8 = shift_i_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_0_9)
      6'b000000 : _zz_shift_q_0_8 = shift_q_map_0;
      6'b000001 : _zz_shift_q_0_8 = shift_q_map_1;
      6'b000010 : _zz_shift_q_0_8 = shift_q_map_2;
      6'b000011 : _zz_shift_q_0_8 = shift_q_map_3;
      6'b000100 : _zz_shift_q_0_8 = shift_q_map_4;
      6'b000101 : _zz_shift_q_0_8 = shift_q_map_5;
      6'b000110 : _zz_shift_q_0_8 = shift_q_map_6;
      6'b000111 : _zz_shift_q_0_8 = shift_q_map_7;
      6'b001000 : _zz_shift_q_0_8 = shift_q_map_8;
      6'b001001 : _zz_shift_q_0_8 = shift_q_map_9;
      6'b001010 : _zz_shift_q_0_8 = shift_q_map_10;
      6'b001011 : _zz_shift_q_0_8 = shift_q_map_11;
      6'b001100 : _zz_shift_q_0_8 = shift_q_map_12;
      6'b001101 : _zz_shift_q_0_8 = shift_q_map_13;
      6'b001110 : _zz_shift_q_0_8 = shift_q_map_14;
      6'b001111 : _zz_shift_q_0_8 = shift_q_map_15;
      6'b010000 : _zz_shift_q_0_8 = shift_q_map_16;
      6'b010001 : _zz_shift_q_0_8 = shift_q_map_17;
      6'b010010 : _zz_shift_q_0_8 = shift_q_map_18;
      6'b010011 : _zz_shift_q_0_8 = shift_q_map_19;
      6'b010100 : _zz_shift_q_0_8 = shift_q_map_20;
      6'b010101 : _zz_shift_q_0_8 = shift_q_map_21;
      6'b010110 : _zz_shift_q_0_8 = shift_q_map_22;
      6'b010111 : _zz_shift_q_0_8 = shift_q_map_23;
      6'b011000 : _zz_shift_q_0_8 = shift_q_map_24;
      6'b011001 : _zz_shift_q_0_8 = shift_q_map_25;
      6'b011010 : _zz_shift_q_0_8 = shift_q_map_26;
      6'b011011 : _zz_shift_q_0_8 = shift_q_map_27;
      6'b011100 : _zz_shift_q_0_8 = shift_q_map_28;
      6'b011101 : _zz_shift_q_0_8 = shift_q_map_29;
      6'b011110 : _zz_shift_q_0_8 = shift_q_map_30;
      6'b011111 : _zz_shift_q_0_8 = shift_q_map_31;
      6'b100000 : _zz_shift_q_0_8 = shift_q_map_32;
      6'b100001 : _zz_shift_q_0_8 = shift_q_map_33;
      6'b100010 : _zz_shift_q_0_8 = shift_q_map_34;
      6'b100011 : _zz_shift_q_0_8 = shift_q_map_35;
      6'b100100 : _zz_shift_q_0_8 = shift_q_map_36;
      6'b100101 : _zz_shift_q_0_8 = shift_q_map_37;
      6'b100110 : _zz_shift_q_0_8 = shift_q_map_38;
      6'b100111 : _zz_shift_q_0_8 = shift_q_map_39;
      6'b101000 : _zz_shift_q_0_8 = shift_q_map_40;
      6'b101001 : _zz_shift_q_0_8 = shift_q_map_41;
      6'b101010 : _zz_shift_q_0_8 = shift_q_map_42;
      6'b101011 : _zz_shift_q_0_8 = shift_q_map_43;
      6'b101100 : _zz_shift_q_0_8 = shift_q_map_44;
      6'b101101 : _zz_shift_q_0_8 = shift_q_map_45;
      6'b101110 : _zz_shift_q_0_8 = shift_q_map_46;
      6'b101111 : _zz_shift_q_0_8 = shift_q_map_47;
      6'b110000 : _zz_shift_q_0_8 = shift_q_map_48;
      6'b110001 : _zz_shift_q_0_8 = shift_q_map_49;
      6'b110010 : _zz_shift_q_0_8 = shift_q_map_50;
      6'b110011 : _zz_shift_q_0_8 = shift_q_map_51;
      6'b110100 : _zz_shift_q_0_8 = shift_q_map_52;
      6'b110101 : _zz_shift_q_0_8 = shift_q_map_53;
      6'b110110 : _zz_shift_q_0_8 = shift_q_map_54;
      6'b110111 : _zz_shift_q_0_8 = shift_q_map_55;
      6'b111000 : _zz_shift_q_0_8 = shift_q_map_56;
      6'b111001 : _zz_shift_q_0_8 = shift_q_map_57;
      6'b111010 : _zz_shift_q_0_8 = shift_q_map_58;
      6'b111011 : _zz_shift_q_0_8 = shift_q_map_59;
      6'b111100 : _zz_shift_q_0_8 = shift_q_map_60;
      6'b111101 : _zz_shift_q_0_8 = shift_q_map_61;
      6'b111110 : _zz_shift_q_0_8 = shift_q_map_62;
      default : _zz_shift_q_0_8 = shift_q_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_1_9)
      6'b000000 : _zz_shift_i_1_8 = shift_i_map_0;
      6'b000001 : _zz_shift_i_1_8 = shift_i_map_1;
      6'b000010 : _zz_shift_i_1_8 = shift_i_map_2;
      6'b000011 : _zz_shift_i_1_8 = shift_i_map_3;
      6'b000100 : _zz_shift_i_1_8 = shift_i_map_4;
      6'b000101 : _zz_shift_i_1_8 = shift_i_map_5;
      6'b000110 : _zz_shift_i_1_8 = shift_i_map_6;
      6'b000111 : _zz_shift_i_1_8 = shift_i_map_7;
      6'b001000 : _zz_shift_i_1_8 = shift_i_map_8;
      6'b001001 : _zz_shift_i_1_8 = shift_i_map_9;
      6'b001010 : _zz_shift_i_1_8 = shift_i_map_10;
      6'b001011 : _zz_shift_i_1_8 = shift_i_map_11;
      6'b001100 : _zz_shift_i_1_8 = shift_i_map_12;
      6'b001101 : _zz_shift_i_1_8 = shift_i_map_13;
      6'b001110 : _zz_shift_i_1_8 = shift_i_map_14;
      6'b001111 : _zz_shift_i_1_8 = shift_i_map_15;
      6'b010000 : _zz_shift_i_1_8 = shift_i_map_16;
      6'b010001 : _zz_shift_i_1_8 = shift_i_map_17;
      6'b010010 : _zz_shift_i_1_8 = shift_i_map_18;
      6'b010011 : _zz_shift_i_1_8 = shift_i_map_19;
      6'b010100 : _zz_shift_i_1_8 = shift_i_map_20;
      6'b010101 : _zz_shift_i_1_8 = shift_i_map_21;
      6'b010110 : _zz_shift_i_1_8 = shift_i_map_22;
      6'b010111 : _zz_shift_i_1_8 = shift_i_map_23;
      6'b011000 : _zz_shift_i_1_8 = shift_i_map_24;
      6'b011001 : _zz_shift_i_1_8 = shift_i_map_25;
      6'b011010 : _zz_shift_i_1_8 = shift_i_map_26;
      6'b011011 : _zz_shift_i_1_8 = shift_i_map_27;
      6'b011100 : _zz_shift_i_1_8 = shift_i_map_28;
      6'b011101 : _zz_shift_i_1_8 = shift_i_map_29;
      6'b011110 : _zz_shift_i_1_8 = shift_i_map_30;
      6'b011111 : _zz_shift_i_1_8 = shift_i_map_31;
      6'b100000 : _zz_shift_i_1_8 = shift_i_map_32;
      6'b100001 : _zz_shift_i_1_8 = shift_i_map_33;
      6'b100010 : _zz_shift_i_1_8 = shift_i_map_34;
      6'b100011 : _zz_shift_i_1_8 = shift_i_map_35;
      6'b100100 : _zz_shift_i_1_8 = shift_i_map_36;
      6'b100101 : _zz_shift_i_1_8 = shift_i_map_37;
      6'b100110 : _zz_shift_i_1_8 = shift_i_map_38;
      6'b100111 : _zz_shift_i_1_8 = shift_i_map_39;
      6'b101000 : _zz_shift_i_1_8 = shift_i_map_40;
      6'b101001 : _zz_shift_i_1_8 = shift_i_map_41;
      6'b101010 : _zz_shift_i_1_8 = shift_i_map_42;
      6'b101011 : _zz_shift_i_1_8 = shift_i_map_43;
      6'b101100 : _zz_shift_i_1_8 = shift_i_map_44;
      6'b101101 : _zz_shift_i_1_8 = shift_i_map_45;
      6'b101110 : _zz_shift_i_1_8 = shift_i_map_46;
      6'b101111 : _zz_shift_i_1_8 = shift_i_map_47;
      6'b110000 : _zz_shift_i_1_8 = shift_i_map_48;
      6'b110001 : _zz_shift_i_1_8 = shift_i_map_49;
      6'b110010 : _zz_shift_i_1_8 = shift_i_map_50;
      6'b110011 : _zz_shift_i_1_8 = shift_i_map_51;
      6'b110100 : _zz_shift_i_1_8 = shift_i_map_52;
      6'b110101 : _zz_shift_i_1_8 = shift_i_map_53;
      6'b110110 : _zz_shift_i_1_8 = shift_i_map_54;
      6'b110111 : _zz_shift_i_1_8 = shift_i_map_55;
      6'b111000 : _zz_shift_i_1_8 = shift_i_map_56;
      6'b111001 : _zz_shift_i_1_8 = shift_i_map_57;
      6'b111010 : _zz_shift_i_1_8 = shift_i_map_58;
      6'b111011 : _zz_shift_i_1_8 = shift_i_map_59;
      6'b111100 : _zz_shift_i_1_8 = shift_i_map_60;
      6'b111101 : _zz_shift_i_1_8 = shift_i_map_61;
      6'b111110 : _zz_shift_i_1_8 = shift_i_map_62;
      default : _zz_shift_i_1_8 = shift_i_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_1_9)
      6'b000000 : _zz_shift_q_1_8 = shift_q_map_0;
      6'b000001 : _zz_shift_q_1_8 = shift_q_map_1;
      6'b000010 : _zz_shift_q_1_8 = shift_q_map_2;
      6'b000011 : _zz_shift_q_1_8 = shift_q_map_3;
      6'b000100 : _zz_shift_q_1_8 = shift_q_map_4;
      6'b000101 : _zz_shift_q_1_8 = shift_q_map_5;
      6'b000110 : _zz_shift_q_1_8 = shift_q_map_6;
      6'b000111 : _zz_shift_q_1_8 = shift_q_map_7;
      6'b001000 : _zz_shift_q_1_8 = shift_q_map_8;
      6'b001001 : _zz_shift_q_1_8 = shift_q_map_9;
      6'b001010 : _zz_shift_q_1_8 = shift_q_map_10;
      6'b001011 : _zz_shift_q_1_8 = shift_q_map_11;
      6'b001100 : _zz_shift_q_1_8 = shift_q_map_12;
      6'b001101 : _zz_shift_q_1_8 = shift_q_map_13;
      6'b001110 : _zz_shift_q_1_8 = shift_q_map_14;
      6'b001111 : _zz_shift_q_1_8 = shift_q_map_15;
      6'b010000 : _zz_shift_q_1_8 = shift_q_map_16;
      6'b010001 : _zz_shift_q_1_8 = shift_q_map_17;
      6'b010010 : _zz_shift_q_1_8 = shift_q_map_18;
      6'b010011 : _zz_shift_q_1_8 = shift_q_map_19;
      6'b010100 : _zz_shift_q_1_8 = shift_q_map_20;
      6'b010101 : _zz_shift_q_1_8 = shift_q_map_21;
      6'b010110 : _zz_shift_q_1_8 = shift_q_map_22;
      6'b010111 : _zz_shift_q_1_8 = shift_q_map_23;
      6'b011000 : _zz_shift_q_1_8 = shift_q_map_24;
      6'b011001 : _zz_shift_q_1_8 = shift_q_map_25;
      6'b011010 : _zz_shift_q_1_8 = shift_q_map_26;
      6'b011011 : _zz_shift_q_1_8 = shift_q_map_27;
      6'b011100 : _zz_shift_q_1_8 = shift_q_map_28;
      6'b011101 : _zz_shift_q_1_8 = shift_q_map_29;
      6'b011110 : _zz_shift_q_1_8 = shift_q_map_30;
      6'b011111 : _zz_shift_q_1_8 = shift_q_map_31;
      6'b100000 : _zz_shift_q_1_8 = shift_q_map_32;
      6'b100001 : _zz_shift_q_1_8 = shift_q_map_33;
      6'b100010 : _zz_shift_q_1_8 = shift_q_map_34;
      6'b100011 : _zz_shift_q_1_8 = shift_q_map_35;
      6'b100100 : _zz_shift_q_1_8 = shift_q_map_36;
      6'b100101 : _zz_shift_q_1_8 = shift_q_map_37;
      6'b100110 : _zz_shift_q_1_8 = shift_q_map_38;
      6'b100111 : _zz_shift_q_1_8 = shift_q_map_39;
      6'b101000 : _zz_shift_q_1_8 = shift_q_map_40;
      6'b101001 : _zz_shift_q_1_8 = shift_q_map_41;
      6'b101010 : _zz_shift_q_1_8 = shift_q_map_42;
      6'b101011 : _zz_shift_q_1_8 = shift_q_map_43;
      6'b101100 : _zz_shift_q_1_8 = shift_q_map_44;
      6'b101101 : _zz_shift_q_1_8 = shift_q_map_45;
      6'b101110 : _zz_shift_q_1_8 = shift_q_map_46;
      6'b101111 : _zz_shift_q_1_8 = shift_q_map_47;
      6'b110000 : _zz_shift_q_1_8 = shift_q_map_48;
      6'b110001 : _zz_shift_q_1_8 = shift_q_map_49;
      6'b110010 : _zz_shift_q_1_8 = shift_q_map_50;
      6'b110011 : _zz_shift_q_1_8 = shift_q_map_51;
      6'b110100 : _zz_shift_q_1_8 = shift_q_map_52;
      6'b110101 : _zz_shift_q_1_8 = shift_q_map_53;
      6'b110110 : _zz_shift_q_1_8 = shift_q_map_54;
      6'b110111 : _zz_shift_q_1_8 = shift_q_map_55;
      6'b111000 : _zz_shift_q_1_8 = shift_q_map_56;
      6'b111001 : _zz_shift_q_1_8 = shift_q_map_57;
      6'b111010 : _zz_shift_q_1_8 = shift_q_map_58;
      6'b111011 : _zz_shift_q_1_8 = shift_q_map_59;
      6'b111100 : _zz_shift_q_1_8 = shift_q_map_60;
      6'b111101 : _zz_shift_q_1_8 = shift_q_map_61;
      6'b111110 : _zz_shift_q_1_8 = shift_q_map_62;
      default : _zz_shift_q_1_8 = shift_q_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_2_9)
      6'b000000 : _zz_shift_i_2_8 = shift_i_map_0;
      6'b000001 : _zz_shift_i_2_8 = shift_i_map_1;
      6'b000010 : _zz_shift_i_2_8 = shift_i_map_2;
      6'b000011 : _zz_shift_i_2_8 = shift_i_map_3;
      6'b000100 : _zz_shift_i_2_8 = shift_i_map_4;
      6'b000101 : _zz_shift_i_2_8 = shift_i_map_5;
      6'b000110 : _zz_shift_i_2_8 = shift_i_map_6;
      6'b000111 : _zz_shift_i_2_8 = shift_i_map_7;
      6'b001000 : _zz_shift_i_2_8 = shift_i_map_8;
      6'b001001 : _zz_shift_i_2_8 = shift_i_map_9;
      6'b001010 : _zz_shift_i_2_8 = shift_i_map_10;
      6'b001011 : _zz_shift_i_2_8 = shift_i_map_11;
      6'b001100 : _zz_shift_i_2_8 = shift_i_map_12;
      6'b001101 : _zz_shift_i_2_8 = shift_i_map_13;
      6'b001110 : _zz_shift_i_2_8 = shift_i_map_14;
      6'b001111 : _zz_shift_i_2_8 = shift_i_map_15;
      6'b010000 : _zz_shift_i_2_8 = shift_i_map_16;
      6'b010001 : _zz_shift_i_2_8 = shift_i_map_17;
      6'b010010 : _zz_shift_i_2_8 = shift_i_map_18;
      6'b010011 : _zz_shift_i_2_8 = shift_i_map_19;
      6'b010100 : _zz_shift_i_2_8 = shift_i_map_20;
      6'b010101 : _zz_shift_i_2_8 = shift_i_map_21;
      6'b010110 : _zz_shift_i_2_8 = shift_i_map_22;
      6'b010111 : _zz_shift_i_2_8 = shift_i_map_23;
      6'b011000 : _zz_shift_i_2_8 = shift_i_map_24;
      6'b011001 : _zz_shift_i_2_8 = shift_i_map_25;
      6'b011010 : _zz_shift_i_2_8 = shift_i_map_26;
      6'b011011 : _zz_shift_i_2_8 = shift_i_map_27;
      6'b011100 : _zz_shift_i_2_8 = shift_i_map_28;
      6'b011101 : _zz_shift_i_2_8 = shift_i_map_29;
      6'b011110 : _zz_shift_i_2_8 = shift_i_map_30;
      6'b011111 : _zz_shift_i_2_8 = shift_i_map_31;
      6'b100000 : _zz_shift_i_2_8 = shift_i_map_32;
      6'b100001 : _zz_shift_i_2_8 = shift_i_map_33;
      6'b100010 : _zz_shift_i_2_8 = shift_i_map_34;
      6'b100011 : _zz_shift_i_2_8 = shift_i_map_35;
      6'b100100 : _zz_shift_i_2_8 = shift_i_map_36;
      6'b100101 : _zz_shift_i_2_8 = shift_i_map_37;
      6'b100110 : _zz_shift_i_2_8 = shift_i_map_38;
      6'b100111 : _zz_shift_i_2_8 = shift_i_map_39;
      6'b101000 : _zz_shift_i_2_8 = shift_i_map_40;
      6'b101001 : _zz_shift_i_2_8 = shift_i_map_41;
      6'b101010 : _zz_shift_i_2_8 = shift_i_map_42;
      6'b101011 : _zz_shift_i_2_8 = shift_i_map_43;
      6'b101100 : _zz_shift_i_2_8 = shift_i_map_44;
      6'b101101 : _zz_shift_i_2_8 = shift_i_map_45;
      6'b101110 : _zz_shift_i_2_8 = shift_i_map_46;
      6'b101111 : _zz_shift_i_2_8 = shift_i_map_47;
      6'b110000 : _zz_shift_i_2_8 = shift_i_map_48;
      6'b110001 : _zz_shift_i_2_8 = shift_i_map_49;
      6'b110010 : _zz_shift_i_2_8 = shift_i_map_50;
      6'b110011 : _zz_shift_i_2_8 = shift_i_map_51;
      6'b110100 : _zz_shift_i_2_8 = shift_i_map_52;
      6'b110101 : _zz_shift_i_2_8 = shift_i_map_53;
      6'b110110 : _zz_shift_i_2_8 = shift_i_map_54;
      6'b110111 : _zz_shift_i_2_8 = shift_i_map_55;
      6'b111000 : _zz_shift_i_2_8 = shift_i_map_56;
      6'b111001 : _zz_shift_i_2_8 = shift_i_map_57;
      6'b111010 : _zz_shift_i_2_8 = shift_i_map_58;
      6'b111011 : _zz_shift_i_2_8 = shift_i_map_59;
      6'b111100 : _zz_shift_i_2_8 = shift_i_map_60;
      6'b111101 : _zz_shift_i_2_8 = shift_i_map_61;
      6'b111110 : _zz_shift_i_2_8 = shift_i_map_62;
      default : _zz_shift_i_2_8 = shift_i_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_2_9)
      6'b000000 : _zz_shift_q_2_8 = shift_q_map_0;
      6'b000001 : _zz_shift_q_2_8 = shift_q_map_1;
      6'b000010 : _zz_shift_q_2_8 = shift_q_map_2;
      6'b000011 : _zz_shift_q_2_8 = shift_q_map_3;
      6'b000100 : _zz_shift_q_2_8 = shift_q_map_4;
      6'b000101 : _zz_shift_q_2_8 = shift_q_map_5;
      6'b000110 : _zz_shift_q_2_8 = shift_q_map_6;
      6'b000111 : _zz_shift_q_2_8 = shift_q_map_7;
      6'b001000 : _zz_shift_q_2_8 = shift_q_map_8;
      6'b001001 : _zz_shift_q_2_8 = shift_q_map_9;
      6'b001010 : _zz_shift_q_2_8 = shift_q_map_10;
      6'b001011 : _zz_shift_q_2_8 = shift_q_map_11;
      6'b001100 : _zz_shift_q_2_8 = shift_q_map_12;
      6'b001101 : _zz_shift_q_2_8 = shift_q_map_13;
      6'b001110 : _zz_shift_q_2_8 = shift_q_map_14;
      6'b001111 : _zz_shift_q_2_8 = shift_q_map_15;
      6'b010000 : _zz_shift_q_2_8 = shift_q_map_16;
      6'b010001 : _zz_shift_q_2_8 = shift_q_map_17;
      6'b010010 : _zz_shift_q_2_8 = shift_q_map_18;
      6'b010011 : _zz_shift_q_2_8 = shift_q_map_19;
      6'b010100 : _zz_shift_q_2_8 = shift_q_map_20;
      6'b010101 : _zz_shift_q_2_8 = shift_q_map_21;
      6'b010110 : _zz_shift_q_2_8 = shift_q_map_22;
      6'b010111 : _zz_shift_q_2_8 = shift_q_map_23;
      6'b011000 : _zz_shift_q_2_8 = shift_q_map_24;
      6'b011001 : _zz_shift_q_2_8 = shift_q_map_25;
      6'b011010 : _zz_shift_q_2_8 = shift_q_map_26;
      6'b011011 : _zz_shift_q_2_8 = shift_q_map_27;
      6'b011100 : _zz_shift_q_2_8 = shift_q_map_28;
      6'b011101 : _zz_shift_q_2_8 = shift_q_map_29;
      6'b011110 : _zz_shift_q_2_8 = shift_q_map_30;
      6'b011111 : _zz_shift_q_2_8 = shift_q_map_31;
      6'b100000 : _zz_shift_q_2_8 = shift_q_map_32;
      6'b100001 : _zz_shift_q_2_8 = shift_q_map_33;
      6'b100010 : _zz_shift_q_2_8 = shift_q_map_34;
      6'b100011 : _zz_shift_q_2_8 = shift_q_map_35;
      6'b100100 : _zz_shift_q_2_8 = shift_q_map_36;
      6'b100101 : _zz_shift_q_2_8 = shift_q_map_37;
      6'b100110 : _zz_shift_q_2_8 = shift_q_map_38;
      6'b100111 : _zz_shift_q_2_8 = shift_q_map_39;
      6'b101000 : _zz_shift_q_2_8 = shift_q_map_40;
      6'b101001 : _zz_shift_q_2_8 = shift_q_map_41;
      6'b101010 : _zz_shift_q_2_8 = shift_q_map_42;
      6'b101011 : _zz_shift_q_2_8 = shift_q_map_43;
      6'b101100 : _zz_shift_q_2_8 = shift_q_map_44;
      6'b101101 : _zz_shift_q_2_8 = shift_q_map_45;
      6'b101110 : _zz_shift_q_2_8 = shift_q_map_46;
      6'b101111 : _zz_shift_q_2_8 = shift_q_map_47;
      6'b110000 : _zz_shift_q_2_8 = shift_q_map_48;
      6'b110001 : _zz_shift_q_2_8 = shift_q_map_49;
      6'b110010 : _zz_shift_q_2_8 = shift_q_map_50;
      6'b110011 : _zz_shift_q_2_8 = shift_q_map_51;
      6'b110100 : _zz_shift_q_2_8 = shift_q_map_52;
      6'b110101 : _zz_shift_q_2_8 = shift_q_map_53;
      6'b110110 : _zz_shift_q_2_8 = shift_q_map_54;
      6'b110111 : _zz_shift_q_2_8 = shift_q_map_55;
      6'b111000 : _zz_shift_q_2_8 = shift_q_map_56;
      6'b111001 : _zz_shift_q_2_8 = shift_q_map_57;
      6'b111010 : _zz_shift_q_2_8 = shift_q_map_58;
      6'b111011 : _zz_shift_q_2_8 = shift_q_map_59;
      6'b111100 : _zz_shift_q_2_8 = shift_q_map_60;
      6'b111101 : _zz_shift_q_2_8 = shift_q_map_61;
      6'b111110 : _zz_shift_q_2_8 = shift_q_map_62;
      default : _zz_shift_q_2_8 = shift_q_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_3_9)
      6'b000000 : _zz_shift_i_3_8 = shift_i_map_0;
      6'b000001 : _zz_shift_i_3_8 = shift_i_map_1;
      6'b000010 : _zz_shift_i_3_8 = shift_i_map_2;
      6'b000011 : _zz_shift_i_3_8 = shift_i_map_3;
      6'b000100 : _zz_shift_i_3_8 = shift_i_map_4;
      6'b000101 : _zz_shift_i_3_8 = shift_i_map_5;
      6'b000110 : _zz_shift_i_3_8 = shift_i_map_6;
      6'b000111 : _zz_shift_i_3_8 = shift_i_map_7;
      6'b001000 : _zz_shift_i_3_8 = shift_i_map_8;
      6'b001001 : _zz_shift_i_3_8 = shift_i_map_9;
      6'b001010 : _zz_shift_i_3_8 = shift_i_map_10;
      6'b001011 : _zz_shift_i_3_8 = shift_i_map_11;
      6'b001100 : _zz_shift_i_3_8 = shift_i_map_12;
      6'b001101 : _zz_shift_i_3_8 = shift_i_map_13;
      6'b001110 : _zz_shift_i_3_8 = shift_i_map_14;
      6'b001111 : _zz_shift_i_3_8 = shift_i_map_15;
      6'b010000 : _zz_shift_i_3_8 = shift_i_map_16;
      6'b010001 : _zz_shift_i_3_8 = shift_i_map_17;
      6'b010010 : _zz_shift_i_3_8 = shift_i_map_18;
      6'b010011 : _zz_shift_i_3_8 = shift_i_map_19;
      6'b010100 : _zz_shift_i_3_8 = shift_i_map_20;
      6'b010101 : _zz_shift_i_3_8 = shift_i_map_21;
      6'b010110 : _zz_shift_i_3_8 = shift_i_map_22;
      6'b010111 : _zz_shift_i_3_8 = shift_i_map_23;
      6'b011000 : _zz_shift_i_3_8 = shift_i_map_24;
      6'b011001 : _zz_shift_i_3_8 = shift_i_map_25;
      6'b011010 : _zz_shift_i_3_8 = shift_i_map_26;
      6'b011011 : _zz_shift_i_3_8 = shift_i_map_27;
      6'b011100 : _zz_shift_i_3_8 = shift_i_map_28;
      6'b011101 : _zz_shift_i_3_8 = shift_i_map_29;
      6'b011110 : _zz_shift_i_3_8 = shift_i_map_30;
      6'b011111 : _zz_shift_i_3_8 = shift_i_map_31;
      6'b100000 : _zz_shift_i_3_8 = shift_i_map_32;
      6'b100001 : _zz_shift_i_3_8 = shift_i_map_33;
      6'b100010 : _zz_shift_i_3_8 = shift_i_map_34;
      6'b100011 : _zz_shift_i_3_8 = shift_i_map_35;
      6'b100100 : _zz_shift_i_3_8 = shift_i_map_36;
      6'b100101 : _zz_shift_i_3_8 = shift_i_map_37;
      6'b100110 : _zz_shift_i_3_8 = shift_i_map_38;
      6'b100111 : _zz_shift_i_3_8 = shift_i_map_39;
      6'b101000 : _zz_shift_i_3_8 = shift_i_map_40;
      6'b101001 : _zz_shift_i_3_8 = shift_i_map_41;
      6'b101010 : _zz_shift_i_3_8 = shift_i_map_42;
      6'b101011 : _zz_shift_i_3_8 = shift_i_map_43;
      6'b101100 : _zz_shift_i_3_8 = shift_i_map_44;
      6'b101101 : _zz_shift_i_3_8 = shift_i_map_45;
      6'b101110 : _zz_shift_i_3_8 = shift_i_map_46;
      6'b101111 : _zz_shift_i_3_8 = shift_i_map_47;
      6'b110000 : _zz_shift_i_3_8 = shift_i_map_48;
      6'b110001 : _zz_shift_i_3_8 = shift_i_map_49;
      6'b110010 : _zz_shift_i_3_8 = shift_i_map_50;
      6'b110011 : _zz_shift_i_3_8 = shift_i_map_51;
      6'b110100 : _zz_shift_i_3_8 = shift_i_map_52;
      6'b110101 : _zz_shift_i_3_8 = shift_i_map_53;
      6'b110110 : _zz_shift_i_3_8 = shift_i_map_54;
      6'b110111 : _zz_shift_i_3_8 = shift_i_map_55;
      6'b111000 : _zz_shift_i_3_8 = shift_i_map_56;
      6'b111001 : _zz_shift_i_3_8 = shift_i_map_57;
      6'b111010 : _zz_shift_i_3_8 = shift_i_map_58;
      6'b111011 : _zz_shift_i_3_8 = shift_i_map_59;
      6'b111100 : _zz_shift_i_3_8 = shift_i_map_60;
      6'b111101 : _zz_shift_i_3_8 = shift_i_map_61;
      6'b111110 : _zz_shift_i_3_8 = shift_i_map_62;
      default : _zz_shift_i_3_8 = shift_i_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_3_9)
      6'b000000 : _zz_shift_q_3_8 = shift_q_map_0;
      6'b000001 : _zz_shift_q_3_8 = shift_q_map_1;
      6'b000010 : _zz_shift_q_3_8 = shift_q_map_2;
      6'b000011 : _zz_shift_q_3_8 = shift_q_map_3;
      6'b000100 : _zz_shift_q_3_8 = shift_q_map_4;
      6'b000101 : _zz_shift_q_3_8 = shift_q_map_5;
      6'b000110 : _zz_shift_q_3_8 = shift_q_map_6;
      6'b000111 : _zz_shift_q_3_8 = shift_q_map_7;
      6'b001000 : _zz_shift_q_3_8 = shift_q_map_8;
      6'b001001 : _zz_shift_q_3_8 = shift_q_map_9;
      6'b001010 : _zz_shift_q_3_8 = shift_q_map_10;
      6'b001011 : _zz_shift_q_3_8 = shift_q_map_11;
      6'b001100 : _zz_shift_q_3_8 = shift_q_map_12;
      6'b001101 : _zz_shift_q_3_8 = shift_q_map_13;
      6'b001110 : _zz_shift_q_3_8 = shift_q_map_14;
      6'b001111 : _zz_shift_q_3_8 = shift_q_map_15;
      6'b010000 : _zz_shift_q_3_8 = shift_q_map_16;
      6'b010001 : _zz_shift_q_3_8 = shift_q_map_17;
      6'b010010 : _zz_shift_q_3_8 = shift_q_map_18;
      6'b010011 : _zz_shift_q_3_8 = shift_q_map_19;
      6'b010100 : _zz_shift_q_3_8 = shift_q_map_20;
      6'b010101 : _zz_shift_q_3_8 = shift_q_map_21;
      6'b010110 : _zz_shift_q_3_8 = shift_q_map_22;
      6'b010111 : _zz_shift_q_3_8 = shift_q_map_23;
      6'b011000 : _zz_shift_q_3_8 = shift_q_map_24;
      6'b011001 : _zz_shift_q_3_8 = shift_q_map_25;
      6'b011010 : _zz_shift_q_3_8 = shift_q_map_26;
      6'b011011 : _zz_shift_q_3_8 = shift_q_map_27;
      6'b011100 : _zz_shift_q_3_8 = shift_q_map_28;
      6'b011101 : _zz_shift_q_3_8 = shift_q_map_29;
      6'b011110 : _zz_shift_q_3_8 = shift_q_map_30;
      6'b011111 : _zz_shift_q_3_8 = shift_q_map_31;
      6'b100000 : _zz_shift_q_3_8 = shift_q_map_32;
      6'b100001 : _zz_shift_q_3_8 = shift_q_map_33;
      6'b100010 : _zz_shift_q_3_8 = shift_q_map_34;
      6'b100011 : _zz_shift_q_3_8 = shift_q_map_35;
      6'b100100 : _zz_shift_q_3_8 = shift_q_map_36;
      6'b100101 : _zz_shift_q_3_8 = shift_q_map_37;
      6'b100110 : _zz_shift_q_3_8 = shift_q_map_38;
      6'b100111 : _zz_shift_q_3_8 = shift_q_map_39;
      6'b101000 : _zz_shift_q_3_8 = shift_q_map_40;
      6'b101001 : _zz_shift_q_3_8 = shift_q_map_41;
      6'b101010 : _zz_shift_q_3_8 = shift_q_map_42;
      6'b101011 : _zz_shift_q_3_8 = shift_q_map_43;
      6'b101100 : _zz_shift_q_3_8 = shift_q_map_44;
      6'b101101 : _zz_shift_q_3_8 = shift_q_map_45;
      6'b101110 : _zz_shift_q_3_8 = shift_q_map_46;
      6'b101111 : _zz_shift_q_3_8 = shift_q_map_47;
      6'b110000 : _zz_shift_q_3_8 = shift_q_map_48;
      6'b110001 : _zz_shift_q_3_8 = shift_q_map_49;
      6'b110010 : _zz_shift_q_3_8 = shift_q_map_50;
      6'b110011 : _zz_shift_q_3_8 = shift_q_map_51;
      6'b110100 : _zz_shift_q_3_8 = shift_q_map_52;
      6'b110101 : _zz_shift_q_3_8 = shift_q_map_53;
      6'b110110 : _zz_shift_q_3_8 = shift_q_map_54;
      6'b110111 : _zz_shift_q_3_8 = shift_q_map_55;
      6'b111000 : _zz_shift_q_3_8 = shift_q_map_56;
      6'b111001 : _zz_shift_q_3_8 = shift_q_map_57;
      6'b111010 : _zz_shift_q_3_8 = shift_q_map_58;
      6'b111011 : _zz_shift_q_3_8 = shift_q_map_59;
      6'b111100 : _zz_shift_q_3_8 = shift_q_map_60;
      6'b111101 : _zz_shift_q_3_8 = shift_q_map_61;
      6'b111110 : _zz_shift_q_3_8 = shift_q_map_62;
      default : _zz_shift_q_3_8 = shift_q_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_4_9)
      6'b000000 : _zz_shift_i_4_8 = shift_i_map_0;
      6'b000001 : _zz_shift_i_4_8 = shift_i_map_1;
      6'b000010 : _zz_shift_i_4_8 = shift_i_map_2;
      6'b000011 : _zz_shift_i_4_8 = shift_i_map_3;
      6'b000100 : _zz_shift_i_4_8 = shift_i_map_4;
      6'b000101 : _zz_shift_i_4_8 = shift_i_map_5;
      6'b000110 : _zz_shift_i_4_8 = shift_i_map_6;
      6'b000111 : _zz_shift_i_4_8 = shift_i_map_7;
      6'b001000 : _zz_shift_i_4_8 = shift_i_map_8;
      6'b001001 : _zz_shift_i_4_8 = shift_i_map_9;
      6'b001010 : _zz_shift_i_4_8 = shift_i_map_10;
      6'b001011 : _zz_shift_i_4_8 = shift_i_map_11;
      6'b001100 : _zz_shift_i_4_8 = shift_i_map_12;
      6'b001101 : _zz_shift_i_4_8 = shift_i_map_13;
      6'b001110 : _zz_shift_i_4_8 = shift_i_map_14;
      6'b001111 : _zz_shift_i_4_8 = shift_i_map_15;
      6'b010000 : _zz_shift_i_4_8 = shift_i_map_16;
      6'b010001 : _zz_shift_i_4_8 = shift_i_map_17;
      6'b010010 : _zz_shift_i_4_8 = shift_i_map_18;
      6'b010011 : _zz_shift_i_4_8 = shift_i_map_19;
      6'b010100 : _zz_shift_i_4_8 = shift_i_map_20;
      6'b010101 : _zz_shift_i_4_8 = shift_i_map_21;
      6'b010110 : _zz_shift_i_4_8 = shift_i_map_22;
      6'b010111 : _zz_shift_i_4_8 = shift_i_map_23;
      6'b011000 : _zz_shift_i_4_8 = shift_i_map_24;
      6'b011001 : _zz_shift_i_4_8 = shift_i_map_25;
      6'b011010 : _zz_shift_i_4_8 = shift_i_map_26;
      6'b011011 : _zz_shift_i_4_8 = shift_i_map_27;
      6'b011100 : _zz_shift_i_4_8 = shift_i_map_28;
      6'b011101 : _zz_shift_i_4_8 = shift_i_map_29;
      6'b011110 : _zz_shift_i_4_8 = shift_i_map_30;
      6'b011111 : _zz_shift_i_4_8 = shift_i_map_31;
      6'b100000 : _zz_shift_i_4_8 = shift_i_map_32;
      6'b100001 : _zz_shift_i_4_8 = shift_i_map_33;
      6'b100010 : _zz_shift_i_4_8 = shift_i_map_34;
      6'b100011 : _zz_shift_i_4_8 = shift_i_map_35;
      6'b100100 : _zz_shift_i_4_8 = shift_i_map_36;
      6'b100101 : _zz_shift_i_4_8 = shift_i_map_37;
      6'b100110 : _zz_shift_i_4_8 = shift_i_map_38;
      6'b100111 : _zz_shift_i_4_8 = shift_i_map_39;
      6'b101000 : _zz_shift_i_4_8 = shift_i_map_40;
      6'b101001 : _zz_shift_i_4_8 = shift_i_map_41;
      6'b101010 : _zz_shift_i_4_8 = shift_i_map_42;
      6'b101011 : _zz_shift_i_4_8 = shift_i_map_43;
      6'b101100 : _zz_shift_i_4_8 = shift_i_map_44;
      6'b101101 : _zz_shift_i_4_8 = shift_i_map_45;
      6'b101110 : _zz_shift_i_4_8 = shift_i_map_46;
      6'b101111 : _zz_shift_i_4_8 = shift_i_map_47;
      6'b110000 : _zz_shift_i_4_8 = shift_i_map_48;
      6'b110001 : _zz_shift_i_4_8 = shift_i_map_49;
      6'b110010 : _zz_shift_i_4_8 = shift_i_map_50;
      6'b110011 : _zz_shift_i_4_8 = shift_i_map_51;
      6'b110100 : _zz_shift_i_4_8 = shift_i_map_52;
      6'b110101 : _zz_shift_i_4_8 = shift_i_map_53;
      6'b110110 : _zz_shift_i_4_8 = shift_i_map_54;
      6'b110111 : _zz_shift_i_4_8 = shift_i_map_55;
      6'b111000 : _zz_shift_i_4_8 = shift_i_map_56;
      6'b111001 : _zz_shift_i_4_8 = shift_i_map_57;
      6'b111010 : _zz_shift_i_4_8 = shift_i_map_58;
      6'b111011 : _zz_shift_i_4_8 = shift_i_map_59;
      6'b111100 : _zz_shift_i_4_8 = shift_i_map_60;
      6'b111101 : _zz_shift_i_4_8 = shift_i_map_61;
      6'b111110 : _zz_shift_i_4_8 = shift_i_map_62;
      default : _zz_shift_i_4_8 = shift_i_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_4_9)
      6'b000000 : _zz_shift_q_4_8 = shift_q_map_0;
      6'b000001 : _zz_shift_q_4_8 = shift_q_map_1;
      6'b000010 : _zz_shift_q_4_8 = shift_q_map_2;
      6'b000011 : _zz_shift_q_4_8 = shift_q_map_3;
      6'b000100 : _zz_shift_q_4_8 = shift_q_map_4;
      6'b000101 : _zz_shift_q_4_8 = shift_q_map_5;
      6'b000110 : _zz_shift_q_4_8 = shift_q_map_6;
      6'b000111 : _zz_shift_q_4_8 = shift_q_map_7;
      6'b001000 : _zz_shift_q_4_8 = shift_q_map_8;
      6'b001001 : _zz_shift_q_4_8 = shift_q_map_9;
      6'b001010 : _zz_shift_q_4_8 = shift_q_map_10;
      6'b001011 : _zz_shift_q_4_8 = shift_q_map_11;
      6'b001100 : _zz_shift_q_4_8 = shift_q_map_12;
      6'b001101 : _zz_shift_q_4_8 = shift_q_map_13;
      6'b001110 : _zz_shift_q_4_8 = shift_q_map_14;
      6'b001111 : _zz_shift_q_4_8 = shift_q_map_15;
      6'b010000 : _zz_shift_q_4_8 = shift_q_map_16;
      6'b010001 : _zz_shift_q_4_8 = shift_q_map_17;
      6'b010010 : _zz_shift_q_4_8 = shift_q_map_18;
      6'b010011 : _zz_shift_q_4_8 = shift_q_map_19;
      6'b010100 : _zz_shift_q_4_8 = shift_q_map_20;
      6'b010101 : _zz_shift_q_4_8 = shift_q_map_21;
      6'b010110 : _zz_shift_q_4_8 = shift_q_map_22;
      6'b010111 : _zz_shift_q_4_8 = shift_q_map_23;
      6'b011000 : _zz_shift_q_4_8 = shift_q_map_24;
      6'b011001 : _zz_shift_q_4_8 = shift_q_map_25;
      6'b011010 : _zz_shift_q_4_8 = shift_q_map_26;
      6'b011011 : _zz_shift_q_4_8 = shift_q_map_27;
      6'b011100 : _zz_shift_q_4_8 = shift_q_map_28;
      6'b011101 : _zz_shift_q_4_8 = shift_q_map_29;
      6'b011110 : _zz_shift_q_4_8 = shift_q_map_30;
      6'b011111 : _zz_shift_q_4_8 = shift_q_map_31;
      6'b100000 : _zz_shift_q_4_8 = shift_q_map_32;
      6'b100001 : _zz_shift_q_4_8 = shift_q_map_33;
      6'b100010 : _zz_shift_q_4_8 = shift_q_map_34;
      6'b100011 : _zz_shift_q_4_8 = shift_q_map_35;
      6'b100100 : _zz_shift_q_4_8 = shift_q_map_36;
      6'b100101 : _zz_shift_q_4_8 = shift_q_map_37;
      6'b100110 : _zz_shift_q_4_8 = shift_q_map_38;
      6'b100111 : _zz_shift_q_4_8 = shift_q_map_39;
      6'b101000 : _zz_shift_q_4_8 = shift_q_map_40;
      6'b101001 : _zz_shift_q_4_8 = shift_q_map_41;
      6'b101010 : _zz_shift_q_4_8 = shift_q_map_42;
      6'b101011 : _zz_shift_q_4_8 = shift_q_map_43;
      6'b101100 : _zz_shift_q_4_8 = shift_q_map_44;
      6'b101101 : _zz_shift_q_4_8 = shift_q_map_45;
      6'b101110 : _zz_shift_q_4_8 = shift_q_map_46;
      6'b101111 : _zz_shift_q_4_8 = shift_q_map_47;
      6'b110000 : _zz_shift_q_4_8 = shift_q_map_48;
      6'b110001 : _zz_shift_q_4_8 = shift_q_map_49;
      6'b110010 : _zz_shift_q_4_8 = shift_q_map_50;
      6'b110011 : _zz_shift_q_4_8 = shift_q_map_51;
      6'b110100 : _zz_shift_q_4_8 = shift_q_map_52;
      6'b110101 : _zz_shift_q_4_8 = shift_q_map_53;
      6'b110110 : _zz_shift_q_4_8 = shift_q_map_54;
      6'b110111 : _zz_shift_q_4_8 = shift_q_map_55;
      6'b111000 : _zz_shift_q_4_8 = shift_q_map_56;
      6'b111001 : _zz_shift_q_4_8 = shift_q_map_57;
      6'b111010 : _zz_shift_q_4_8 = shift_q_map_58;
      6'b111011 : _zz_shift_q_4_8 = shift_q_map_59;
      6'b111100 : _zz_shift_q_4_8 = shift_q_map_60;
      6'b111101 : _zz_shift_q_4_8 = shift_q_map_61;
      6'b111110 : _zz_shift_q_4_8 = shift_q_map_62;
      default : _zz_shift_q_4_8 = shift_q_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_5_9)
      6'b000000 : _zz_shift_i_5_8 = shift_i_map_0;
      6'b000001 : _zz_shift_i_5_8 = shift_i_map_1;
      6'b000010 : _zz_shift_i_5_8 = shift_i_map_2;
      6'b000011 : _zz_shift_i_5_8 = shift_i_map_3;
      6'b000100 : _zz_shift_i_5_8 = shift_i_map_4;
      6'b000101 : _zz_shift_i_5_8 = shift_i_map_5;
      6'b000110 : _zz_shift_i_5_8 = shift_i_map_6;
      6'b000111 : _zz_shift_i_5_8 = shift_i_map_7;
      6'b001000 : _zz_shift_i_5_8 = shift_i_map_8;
      6'b001001 : _zz_shift_i_5_8 = shift_i_map_9;
      6'b001010 : _zz_shift_i_5_8 = shift_i_map_10;
      6'b001011 : _zz_shift_i_5_8 = shift_i_map_11;
      6'b001100 : _zz_shift_i_5_8 = shift_i_map_12;
      6'b001101 : _zz_shift_i_5_8 = shift_i_map_13;
      6'b001110 : _zz_shift_i_5_8 = shift_i_map_14;
      6'b001111 : _zz_shift_i_5_8 = shift_i_map_15;
      6'b010000 : _zz_shift_i_5_8 = shift_i_map_16;
      6'b010001 : _zz_shift_i_5_8 = shift_i_map_17;
      6'b010010 : _zz_shift_i_5_8 = shift_i_map_18;
      6'b010011 : _zz_shift_i_5_8 = shift_i_map_19;
      6'b010100 : _zz_shift_i_5_8 = shift_i_map_20;
      6'b010101 : _zz_shift_i_5_8 = shift_i_map_21;
      6'b010110 : _zz_shift_i_5_8 = shift_i_map_22;
      6'b010111 : _zz_shift_i_5_8 = shift_i_map_23;
      6'b011000 : _zz_shift_i_5_8 = shift_i_map_24;
      6'b011001 : _zz_shift_i_5_8 = shift_i_map_25;
      6'b011010 : _zz_shift_i_5_8 = shift_i_map_26;
      6'b011011 : _zz_shift_i_5_8 = shift_i_map_27;
      6'b011100 : _zz_shift_i_5_8 = shift_i_map_28;
      6'b011101 : _zz_shift_i_5_8 = shift_i_map_29;
      6'b011110 : _zz_shift_i_5_8 = shift_i_map_30;
      6'b011111 : _zz_shift_i_5_8 = shift_i_map_31;
      6'b100000 : _zz_shift_i_5_8 = shift_i_map_32;
      6'b100001 : _zz_shift_i_5_8 = shift_i_map_33;
      6'b100010 : _zz_shift_i_5_8 = shift_i_map_34;
      6'b100011 : _zz_shift_i_5_8 = shift_i_map_35;
      6'b100100 : _zz_shift_i_5_8 = shift_i_map_36;
      6'b100101 : _zz_shift_i_5_8 = shift_i_map_37;
      6'b100110 : _zz_shift_i_5_8 = shift_i_map_38;
      6'b100111 : _zz_shift_i_5_8 = shift_i_map_39;
      6'b101000 : _zz_shift_i_5_8 = shift_i_map_40;
      6'b101001 : _zz_shift_i_5_8 = shift_i_map_41;
      6'b101010 : _zz_shift_i_5_8 = shift_i_map_42;
      6'b101011 : _zz_shift_i_5_8 = shift_i_map_43;
      6'b101100 : _zz_shift_i_5_8 = shift_i_map_44;
      6'b101101 : _zz_shift_i_5_8 = shift_i_map_45;
      6'b101110 : _zz_shift_i_5_8 = shift_i_map_46;
      6'b101111 : _zz_shift_i_5_8 = shift_i_map_47;
      6'b110000 : _zz_shift_i_5_8 = shift_i_map_48;
      6'b110001 : _zz_shift_i_5_8 = shift_i_map_49;
      6'b110010 : _zz_shift_i_5_8 = shift_i_map_50;
      6'b110011 : _zz_shift_i_5_8 = shift_i_map_51;
      6'b110100 : _zz_shift_i_5_8 = shift_i_map_52;
      6'b110101 : _zz_shift_i_5_8 = shift_i_map_53;
      6'b110110 : _zz_shift_i_5_8 = shift_i_map_54;
      6'b110111 : _zz_shift_i_5_8 = shift_i_map_55;
      6'b111000 : _zz_shift_i_5_8 = shift_i_map_56;
      6'b111001 : _zz_shift_i_5_8 = shift_i_map_57;
      6'b111010 : _zz_shift_i_5_8 = shift_i_map_58;
      6'b111011 : _zz_shift_i_5_8 = shift_i_map_59;
      6'b111100 : _zz_shift_i_5_8 = shift_i_map_60;
      6'b111101 : _zz_shift_i_5_8 = shift_i_map_61;
      6'b111110 : _zz_shift_i_5_8 = shift_i_map_62;
      default : _zz_shift_i_5_8 = shift_i_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_5_9)
      6'b000000 : _zz_shift_q_5_8 = shift_q_map_0;
      6'b000001 : _zz_shift_q_5_8 = shift_q_map_1;
      6'b000010 : _zz_shift_q_5_8 = shift_q_map_2;
      6'b000011 : _zz_shift_q_5_8 = shift_q_map_3;
      6'b000100 : _zz_shift_q_5_8 = shift_q_map_4;
      6'b000101 : _zz_shift_q_5_8 = shift_q_map_5;
      6'b000110 : _zz_shift_q_5_8 = shift_q_map_6;
      6'b000111 : _zz_shift_q_5_8 = shift_q_map_7;
      6'b001000 : _zz_shift_q_5_8 = shift_q_map_8;
      6'b001001 : _zz_shift_q_5_8 = shift_q_map_9;
      6'b001010 : _zz_shift_q_5_8 = shift_q_map_10;
      6'b001011 : _zz_shift_q_5_8 = shift_q_map_11;
      6'b001100 : _zz_shift_q_5_8 = shift_q_map_12;
      6'b001101 : _zz_shift_q_5_8 = shift_q_map_13;
      6'b001110 : _zz_shift_q_5_8 = shift_q_map_14;
      6'b001111 : _zz_shift_q_5_8 = shift_q_map_15;
      6'b010000 : _zz_shift_q_5_8 = shift_q_map_16;
      6'b010001 : _zz_shift_q_5_8 = shift_q_map_17;
      6'b010010 : _zz_shift_q_5_8 = shift_q_map_18;
      6'b010011 : _zz_shift_q_5_8 = shift_q_map_19;
      6'b010100 : _zz_shift_q_5_8 = shift_q_map_20;
      6'b010101 : _zz_shift_q_5_8 = shift_q_map_21;
      6'b010110 : _zz_shift_q_5_8 = shift_q_map_22;
      6'b010111 : _zz_shift_q_5_8 = shift_q_map_23;
      6'b011000 : _zz_shift_q_5_8 = shift_q_map_24;
      6'b011001 : _zz_shift_q_5_8 = shift_q_map_25;
      6'b011010 : _zz_shift_q_5_8 = shift_q_map_26;
      6'b011011 : _zz_shift_q_5_8 = shift_q_map_27;
      6'b011100 : _zz_shift_q_5_8 = shift_q_map_28;
      6'b011101 : _zz_shift_q_5_8 = shift_q_map_29;
      6'b011110 : _zz_shift_q_5_8 = shift_q_map_30;
      6'b011111 : _zz_shift_q_5_8 = shift_q_map_31;
      6'b100000 : _zz_shift_q_5_8 = shift_q_map_32;
      6'b100001 : _zz_shift_q_5_8 = shift_q_map_33;
      6'b100010 : _zz_shift_q_5_8 = shift_q_map_34;
      6'b100011 : _zz_shift_q_5_8 = shift_q_map_35;
      6'b100100 : _zz_shift_q_5_8 = shift_q_map_36;
      6'b100101 : _zz_shift_q_5_8 = shift_q_map_37;
      6'b100110 : _zz_shift_q_5_8 = shift_q_map_38;
      6'b100111 : _zz_shift_q_5_8 = shift_q_map_39;
      6'b101000 : _zz_shift_q_5_8 = shift_q_map_40;
      6'b101001 : _zz_shift_q_5_8 = shift_q_map_41;
      6'b101010 : _zz_shift_q_5_8 = shift_q_map_42;
      6'b101011 : _zz_shift_q_5_8 = shift_q_map_43;
      6'b101100 : _zz_shift_q_5_8 = shift_q_map_44;
      6'b101101 : _zz_shift_q_5_8 = shift_q_map_45;
      6'b101110 : _zz_shift_q_5_8 = shift_q_map_46;
      6'b101111 : _zz_shift_q_5_8 = shift_q_map_47;
      6'b110000 : _zz_shift_q_5_8 = shift_q_map_48;
      6'b110001 : _zz_shift_q_5_8 = shift_q_map_49;
      6'b110010 : _zz_shift_q_5_8 = shift_q_map_50;
      6'b110011 : _zz_shift_q_5_8 = shift_q_map_51;
      6'b110100 : _zz_shift_q_5_8 = shift_q_map_52;
      6'b110101 : _zz_shift_q_5_8 = shift_q_map_53;
      6'b110110 : _zz_shift_q_5_8 = shift_q_map_54;
      6'b110111 : _zz_shift_q_5_8 = shift_q_map_55;
      6'b111000 : _zz_shift_q_5_8 = shift_q_map_56;
      6'b111001 : _zz_shift_q_5_8 = shift_q_map_57;
      6'b111010 : _zz_shift_q_5_8 = shift_q_map_58;
      6'b111011 : _zz_shift_q_5_8 = shift_q_map_59;
      6'b111100 : _zz_shift_q_5_8 = shift_q_map_60;
      6'b111101 : _zz_shift_q_5_8 = shift_q_map_61;
      6'b111110 : _zz_shift_q_5_8 = shift_q_map_62;
      default : _zz_shift_q_5_8 = shift_q_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_6_9)
      6'b000000 : _zz_shift_i_6_8 = shift_i_map_0;
      6'b000001 : _zz_shift_i_6_8 = shift_i_map_1;
      6'b000010 : _zz_shift_i_6_8 = shift_i_map_2;
      6'b000011 : _zz_shift_i_6_8 = shift_i_map_3;
      6'b000100 : _zz_shift_i_6_8 = shift_i_map_4;
      6'b000101 : _zz_shift_i_6_8 = shift_i_map_5;
      6'b000110 : _zz_shift_i_6_8 = shift_i_map_6;
      6'b000111 : _zz_shift_i_6_8 = shift_i_map_7;
      6'b001000 : _zz_shift_i_6_8 = shift_i_map_8;
      6'b001001 : _zz_shift_i_6_8 = shift_i_map_9;
      6'b001010 : _zz_shift_i_6_8 = shift_i_map_10;
      6'b001011 : _zz_shift_i_6_8 = shift_i_map_11;
      6'b001100 : _zz_shift_i_6_8 = shift_i_map_12;
      6'b001101 : _zz_shift_i_6_8 = shift_i_map_13;
      6'b001110 : _zz_shift_i_6_8 = shift_i_map_14;
      6'b001111 : _zz_shift_i_6_8 = shift_i_map_15;
      6'b010000 : _zz_shift_i_6_8 = shift_i_map_16;
      6'b010001 : _zz_shift_i_6_8 = shift_i_map_17;
      6'b010010 : _zz_shift_i_6_8 = shift_i_map_18;
      6'b010011 : _zz_shift_i_6_8 = shift_i_map_19;
      6'b010100 : _zz_shift_i_6_8 = shift_i_map_20;
      6'b010101 : _zz_shift_i_6_8 = shift_i_map_21;
      6'b010110 : _zz_shift_i_6_8 = shift_i_map_22;
      6'b010111 : _zz_shift_i_6_8 = shift_i_map_23;
      6'b011000 : _zz_shift_i_6_8 = shift_i_map_24;
      6'b011001 : _zz_shift_i_6_8 = shift_i_map_25;
      6'b011010 : _zz_shift_i_6_8 = shift_i_map_26;
      6'b011011 : _zz_shift_i_6_8 = shift_i_map_27;
      6'b011100 : _zz_shift_i_6_8 = shift_i_map_28;
      6'b011101 : _zz_shift_i_6_8 = shift_i_map_29;
      6'b011110 : _zz_shift_i_6_8 = shift_i_map_30;
      6'b011111 : _zz_shift_i_6_8 = shift_i_map_31;
      6'b100000 : _zz_shift_i_6_8 = shift_i_map_32;
      6'b100001 : _zz_shift_i_6_8 = shift_i_map_33;
      6'b100010 : _zz_shift_i_6_8 = shift_i_map_34;
      6'b100011 : _zz_shift_i_6_8 = shift_i_map_35;
      6'b100100 : _zz_shift_i_6_8 = shift_i_map_36;
      6'b100101 : _zz_shift_i_6_8 = shift_i_map_37;
      6'b100110 : _zz_shift_i_6_8 = shift_i_map_38;
      6'b100111 : _zz_shift_i_6_8 = shift_i_map_39;
      6'b101000 : _zz_shift_i_6_8 = shift_i_map_40;
      6'b101001 : _zz_shift_i_6_8 = shift_i_map_41;
      6'b101010 : _zz_shift_i_6_8 = shift_i_map_42;
      6'b101011 : _zz_shift_i_6_8 = shift_i_map_43;
      6'b101100 : _zz_shift_i_6_8 = shift_i_map_44;
      6'b101101 : _zz_shift_i_6_8 = shift_i_map_45;
      6'b101110 : _zz_shift_i_6_8 = shift_i_map_46;
      6'b101111 : _zz_shift_i_6_8 = shift_i_map_47;
      6'b110000 : _zz_shift_i_6_8 = shift_i_map_48;
      6'b110001 : _zz_shift_i_6_8 = shift_i_map_49;
      6'b110010 : _zz_shift_i_6_8 = shift_i_map_50;
      6'b110011 : _zz_shift_i_6_8 = shift_i_map_51;
      6'b110100 : _zz_shift_i_6_8 = shift_i_map_52;
      6'b110101 : _zz_shift_i_6_8 = shift_i_map_53;
      6'b110110 : _zz_shift_i_6_8 = shift_i_map_54;
      6'b110111 : _zz_shift_i_6_8 = shift_i_map_55;
      6'b111000 : _zz_shift_i_6_8 = shift_i_map_56;
      6'b111001 : _zz_shift_i_6_8 = shift_i_map_57;
      6'b111010 : _zz_shift_i_6_8 = shift_i_map_58;
      6'b111011 : _zz_shift_i_6_8 = shift_i_map_59;
      6'b111100 : _zz_shift_i_6_8 = shift_i_map_60;
      6'b111101 : _zz_shift_i_6_8 = shift_i_map_61;
      6'b111110 : _zz_shift_i_6_8 = shift_i_map_62;
      default : _zz_shift_i_6_8 = shift_i_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_6_9)
      6'b000000 : _zz_shift_q_6_8 = shift_q_map_0;
      6'b000001 : _zz_shift_q_6_8 = shift_q_map_1;
      6'b000010 : _zz_shift_q_6_8 = shift_q_map_2;
      6'b000011 : _zz_shift_q_6_8 = shift_q_map_3;
      6'b000100 : _zz_shift_q_6_8 = shift_q_map_4;
      6'b000101 : _zz_shift_q_6_8 = shift_q_map_5;
      6'b000110 : _zz_shift_q_6_8 = shift_q_map_6;
      6'b000111 : _zz_shift_q_6_8 = shift_q_map_7;
      6'b001000 : _zz_shift_q_6_8 = shift_q_map_8;
      6'b001001 : _zz_shift_q_6_8 = shift_q_map_9;
      6'b001010 : _zz_shift_q_6_8 = shift_q_map_10;
      6'b001011 : _zz_shift_q_6_8 = shift_q_map_11;
      6'b001100 : _zz_shift_q_6_8 = shift_q_map_12;
      6'b001101 : _zz_shift_q_6_8 = shift_q_map_13;
      6'b001110 : _zz_shift_q_6_8 = shift_q_map_14;
      6'b001111 : _zz_shift_q_6_8 = shift_q_map_15;
      6'b010000 : _zz_shift_q_6_8 = shift_q_map_16;
      6'b010001 : _zz_shift_q_6_8 = shift_q_map_17;
      6'b010010 : _zz_shift_q_6_8 = shift_q_map_18;
      6'b010011 : _zz_shift_q_6_8 = shift_q_map_19;
      6'b010100 : _zz_shift_q_6_8 = shift_q_map_20;
      6'b010101 : _zz_shift_q_6_8 = shift_q_map_21;
      6'b010110 : _zz_shift_q_6_8 = shift_q_map_22;
      6'b010111 : _zz_shift_q_6_8 = shift_q_map_23;
      6'b011000 : _zz_shift_q_6_8 = shift_q_map_24;
      6'b011001 : _zz_shift_q_6_8 = shift_q_map_25;
      6'b011010 : _zz_shift_q_6_8 = shift_q_map_26;
      6'b011011 : _zz_shift_q_6_8 = shift_q_map_27;
      6'b011100 : _zz_shift_q_6_8 = shift_q_map_28;
      6'b011101 : _zz_shift_q_6_8 = shift_q_map_29;
      6'b011110 : _zz_shift_q_6_8 = shift_q_map_30;
      6'b011111 : _zz_shift_q_6_8 = shift_q_map_31;
      6'b100000 : _zz_shift_q_6_8 = shift_q_map_32;
      6'b100001 : _zz_shift_q_6_8 = shift_q_map_33;
      6'b100010 : _zz_shift_q_6_8 = shift_q_map_34;
      6'b100011 : _zz_shift_q_6_8 = shift_q_map_35;
      6'b100100 : _zz_shift_q_6_8 = shift_q_map_36;
      6'b100101 : _zz_shift_q_6_8 = shift_q_map_37;
      6'b100110 : _zz_shift_q_6_8 = shift_q_map_38;
      6'b100111 : _zz_shift_q_6_8 = shift_q_map_39;
      6'b101000 : _zz_shift_q_6_8 = shift_q_map_40;
      6'b101001 : _zz_shift_q_6_8 = shift_q_map_41;
      6'b101010 : _zz_shift_q_6_8 = shift_q_map_42;
      6'b101011 : _zz_shift_q_6_8 = shift_q_map_43;
      6'b101100 : _zz_shift_q_6_8 = shift_q_map_44;
      6'b101101 : _zz_shift_q_6_8 = shift_q_map_45;
      6'b101110 : _zz_shift_q_6_8 = shift_q_map_46;
      6'b101111 : _zz_shift_q_6_8 = shift_q_map_47;
      6'b110000 : _zz_shift_q_6_8 = shift_q_map_48;
      6'b110001 : _zz_shift_q_6_8 = shift_q_map_49;
      6'b110010 : _zz_shift_q_6_8 = shift_q_map_50;
      6'b110011 : _zz_shift_q_6_8 = shift_q_map_51;
      6'b110100 : _zz_shift_q_6_8 = shift_q_map_52;
      6'b110101 : _zz_shift_q_6_8 = shift_q_map_53;
      6'b110110 : _zz_shift_q_6_8 = shift_q_map_54;
      6'b110111 : _zz_shift_q_6_8 = shift_q_map_55;
      6'b111000 : _zz_shift_q_6_8 = shift_q_map_56;
      6'b111001 : _zz_shift_q_6_8 = shift_q_map_57;
      6'b111010 : _zz_shift_q_6_8 = shift_q_map_58;
      6'b111011 : _zz_shift_q_6_8 = shift_q_map_59;
      6'b111100 : _zz_shift_q_6_8 = shift_q_map_60;
      6'b111101 : _zz_shift_q_6_8 = shift_q_map_61;
      6'b111110 : _zz_shift_q_6_8 = shift_q_map_62;
      default : _zz_shift_q_6_8 = shift_q_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_7_9)
      6'b000000 : _zz_shift_i_7_8 = shift_i_map_0;
      6'b000001 : _zz_shift_i_7_8 = shift_i_map_1;
      6'b000010 : _zz_shift_i_7_8 = shift_i_map_2;
      6'b000011 : _zz_shift_i_7_8 = shift_i_map_3;
      6'b000100 : _zz_shift_i_7_8 = shift_i_map_4;
      6'b000101 : _zz_shift_i_7_8 = shift_i_map_5;
      6'b000110 : _zz_shift_i_7_8 = shift_i_map_6;
      6'b000111 : _zz_shift_i_7_8 = shift_i_map_7;
      6'b001000 : _zz_shift_i_7_8 = shift_i_map_8;
      6'b001001 : _zz_shift_i_7_8 = shift_i_map_9;
      6'b001010 : _zz_shift_i_7_8 = shift_i_map_10;
      6'b001011 : _zz_shift_i_7_8 = shift_i_map_11;
      6'b001100 : _zz_shift_i_7_8 = shift_i_map_12;
      6'b001101 : _zz_shift_i_7_8 = shift_i_map_13;
      6'b001110 : _zz_shift_i_7_8 = shift_i_map_14;
      6'b001111 : _zz_shift_i_7_8 = shift_i_map_15;
      6'b010000 : _zz_shift_i_7_8 = shift_i_map_16;
      6'b010001 : _zz_shift_i_7_8 = shift_i_map_17;
      6'b010010 : _zz_shift_i_7_8 = shift_i_map_18;
      6'b010011 : _zz_shift_i_7_8 = shift_i_map_19;
      6'b010100 : _zz_shift_i_7_8 = shift_i_map_20;
      6'b010101 : _zz_shift_i_7_8 = shift_i_map_21;
      6'b010110 : _zz_shift_i_7_8 = shift_i_map_22;
      6'b010111 : _zz_shift_i_7_8 = shift_i_map_23;
      6'b011000 : _zz_shift_i_7_8 = shift_i_map_24;
      6'b011001 : _zz_shift_i_7_8 = shift_i_map_25;
      6'b011010 : _zz_shift_i_7_8 = shift_i_map_26;
      6'b011011 : _zz_shift_i_7_8 = shift_i_map_27;
      6'b011100 : _zz_shift_i_7_8 = shift_i_map_28;
      6'b011101 : _zz_shift_i_7_8 = shift_i_map_29;
      6'b011110 : _zz_shift_i_7_8 = shift_i_map_30;
      6'b011111 : _zz_shift_i_7_8 = shift_i_map_31;
      6'b100000 : _zz_shift_i_7_8 = shift_i_map_32;
      6'b100001 : _zz_shift_i_7_8 = shift_i_map_33;
      6'b100010 : _zz_shift_i_7_8 = shift_i_map_34;
      6'b100011 : _zz_shift_i_7_8 = shift_i_map_35;
      6'b100100 : _zz_shift_i_7_8 = shift_i_map_36;
      6'b100101 : _zz_shift_i_7_8 = shift_i_map_37;
      6'b100110 : _zz_shift_i_7_8 = shift_i_map_38;
      6'b100111 : _zz_shift_i_7_8 = shift_i_map_39;
      6'b101000 : _zz_shift_i_7_8 = shift_i_map_40;
      6'b101001 : _zz_shift_i_7_8 = shift_i_map_41;
      6'b101010 : _zz_shift_i_7_8 = shift_i_map_42;
      6'b101011 : _zz_shift_i_7_8 = shift_i_map_43;
      6'b101100 : _zz_shift_i_7_8 = shift_i_map_44;
      6'b101101 : _zz_shift_i_7_8 = shift_i_map_45;
      6'b101110 : _zz_shift_i_7_8 = shift_i_map_46;
      6'b101111 : _zz_shift_i_7_8 = shift_i_map_47;
      6'b110000 : _zz_shift_i_7_8 = shift_i_map_48;
      6'b110001 : _zz_shift_i_7_8 = shift_i_map_49;
      6'b110010 : _zz_shift_i_7_8 = shift_i_map_50;
      6'b110011 : _zz_shift_i_7_8 = shift_i_map_51;
      6'b110100 : _zz_shift_i_7_8 = shift_i_map_52;
      6'b110101 : _zz_shift_i_7_8 = shift_i_map_53;
      6'b110110 : _zz_shift_i_7_8 = shift_i_map_54;
      6'b110111 : _zz_shift_i_7_8 = shift_i_map_55;
      6'b111000 : _zz_shift_i_7_8 = shift_i_map_56;
      6'b111001 : _zz_shift_i_7_8 = shift_i_map_57;
      6'b111010 : _zz_shift_i_7_8 = shift_i_map_58;
      6'b111011 : _zz_shift_i_7_8 = shift_i_map_59;
      6'b111100 : _zz_shift_i_7_8 = shift_i_map_60;
      6'b111101 : _zz_shift_i_7_8 = shift_i_map_61;
      6'b111110 : _zz_shift_i_7_8 = shift_i_map_62;
      default : _zz_shift_i_7_8 = shift_i_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_7_9)
      6'b000000 : _zz_shift_q_7_8 = shift_q_map_0;
      6'b000001 : _zz_shift_q_7_8 = shift_q_map_1;
      6'b000010 : _zz_shift_q_7_8 = shift_q_map_2;
      6'b000011 : _zz_shift_q_7_8 = shift_q_map_3;
      6'b000100 : _zz_shift_q_7_8 = shift_q_map_4;
      6'b000101 : _zz_shift_q_7_8 = shift_q_map_5;
      6'b000110 : _zz_shift_q_7_8 = shift_q_map_6;
      6'b000111 : _zz_shift_q_7_8 = shift_q_map_7;
      6'b001000 : _zz_shift_q_7_8 = shift_q_map_8;
      6'b001001 : _zz_shift_q_7_8 = shift_q_map_9;
      6'b001010 : _zz_shift_q_7_8 = shift_q_map_10;
      6'b001011 : _zz_shift_q_7_8 = shift_q_map_11;
      6'b001100 : _zz_shift_q_7_8 = shift_q_map_12;
      6'b001101 : _zz_shift_q_7_8 = shift_q_map_13;
      6'b001110 : _zz_shift_q_7_8 = shift_q_map_14;
      6'b001111 : _zz_shift_q_7_8 = shift_q_map_15;
      6'b010000 : _zz_shift_q_7_8 = shift_q_map_16;
      6'b010001 : _zz_shift_q_7_8 = shift_q_map_17;
      6'b010010 : _zz_shift_q_7_8 = shift_q_map_18;
      6'b010011 : _zz_shift_q_7_8 = shift_q_map_19;
      6'b010100 : _zz_shift_q_7_8 = shift_q_map_20;
      6'b010101 : _zz_shift_q_7_8 = shift_q_map_21;
      6'b010110 : _zz_shift_q_7_8 = shift_q_map_22;
      6'b010111 : _zz_shift_q_7_8 = shift_q_map_23;
      6'b011000 : _zz_shift_q_7_8 = shift_q_map_24;
      6'b011001 : _zz_shift_q_7_8 = shift_q_map_25;
      6'b011010 : _zz_shift_q_7_8 = shift_q_map_26;
      6'b011011 : _zz_shift_q_7_8 = shift_q_map_27;
      6'b011100 : _zz_shift_q_7_8 = shift_q_map_28;
      6'b011101 : _zz_shift_q_7_8 = shift_q_map_29;
      6'b011110 : _zz_shift_q_7_8 = shift_q_map_30;
      6'b011111 : _zz_shift_q_7_8 = shift_q_map_31;
      6'b100000 : _zz_shift_q_7_8 = shift_q_map_32;
      6'b100001 : _zz_shift_q_7_8 = shift_q_map_33;
      6'b100010 : _zz_shift_q_7_8 = shift_q_map_34;
      6'b100011 : _zz_shift_q_7_8 = shift_q_map_35;
      6'b100100 : _zz_shift_q_7_8 = shift_q_map_36;
      6'b100101 : _zz_shift_q_7_8 = shift_q_map_37;
      6'b100110 : _zz_shift_q_7_8 = shift_q_map_38;
      6'b100111 : _zz_shift_q_7_8 = shift_q_map_39;
      6'b101000 : _zz_shift_q_7_8 = shift_q_map_40;
      6'b101001 : _zz_shift_q_7_8 = shift_q_map_41;
      6'b101010 : _zz_shift_q_7_8 = shift_q_map_42;
      6'b101011 : _zz_shift_q_7_8 = shift_q_map_43;
      6'b101100 : _zz_shift_q_7_8 = shift_q_map_44;
      6'b101101 : _zz_shift_q_7_8 = shift_q_map_45;
      6'b101110 : _zz_shift_q_7_8 = shift_q_map_46;
      6'b101111 : _zz_shift_q_7_8 = shift_q_map_47;
      6'b110000 : _zz_shift_q_7_8 = shift_q_map_48;
      6'b110001 : _zz_shift_q_7_8 = shift_q_map_49;
      6'b110010 : _zz_shift_q_7_8 = shift_q_map_50;
      6'b110011 : _zz_shift_q_7_8 = shift_q_map_51;
      6'b110100 : _zz_shift_q_7_8 = shift_q_map_52;
      6'b110101 : _zz_shift_q_7_8 = shift_q_map_53;
      6'b110110 : _zz_shift_q_7_8 = shift_q_map_54;
      6'b110111 : _zz_shift_q_7_8 = shift_q_map_55;
      6'b111000 : _zz_shift_q_7_8 = shift_q_map_56;
      6'b111001 : _zz_shift_q_7_8 = shift_q_map_57;
      6'b111010 : _zz_shift_q_7_8 = shift_q_map_58;
      6'b111011 : _zz_shift_q_7_8 = shift_q_map_59;
      6'b111100 : _zz_shift_q_7_8 = shift_q_map_60;
      6'b111101 : _zz_shift_q_7_8 = shift_q_map_61;
      6'b111110 : _zz_shift_q_7_8 = shift_q_map_62;
      default : _zz_shift_q_7_8 = shift_q_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_0_11)
      6'b000000 : _zz_shift_i_0_10 = shift_i_map_0;
      6'b000001 : _zz_shift_i_0_10 = shift_i_map_1;
      6'b000010 : _zz_shift_i_0_10 = shift_i_map_2;
      6'b000011 : _zz_shift_i_0_10 = shift_i_map_3;
      6'b000100 : _zz_shift_i_0_10 = shift_i_map_4;
      6'b000101 : _zz_shift_i_0_10 = shift_i_map_5;
      6'b000110 : _zz_shift_i_0_10 = shift_i_map_6;
      6'b000111 : _zz_shift_i_0_10 = shift_i_map_7;
      6'b001000 : _zz_shift_i_0_10 = shift_i_map_8;
      6'b001001 : _zz_shift_i_0_10 = shift_i_map_9;
      6'b001010 : _zz_shift_i_0_10 = shift_i_map_10;
      6'b001011 : _zz_shift_i_0_10 = shift_i_map_11;
      6'b001100 : _zz_shift_i_0_10 = shift_i_map_12;
      6'b001101 : _zz_shift_i_0_10 = shift_i_map_13;
      6'b001110 : _zz_shift_i_0_10 = shift_i_map_14;
      6'b001111 : _zz_shift_i_0_10 = shift_i_map_15;
      6'b010000 : _zz_shift_i_0_10 = shift_i_map_16;
      6'b010001 : _zz_shift_i_0_10 = shift_i_map_17;
      6'b010010 : _zz_shift_i_0_10 = shift_i_map_18;
      6'b010011 : _zz_shift_i_0_10 = shift_i_map_19;
      6'b010100 : _zz_shift_i_0_10 = shift_i_map_20;
      6'b010101 : _zz_shift_i_0_10 = shift_i_map_21;
      6'b010110 : _zz_shift_i_0_10 = shift_i_map_22;
      6'b010111 : _zz_shift_i_0_10 = shift_i_map_23;
      6'b011000 : _zz_shift_i_0_10 = shift_i_map_24;
      6'b011001 : _zz_shift_i_0_10 = shift_i_map_25;
      6'b011010 : _zz_shift_i_0_10 = shift_i_map_26;
      6'b011011 : _zz_shift_i_0_10 = shift_i_map_27;
      6'b011100 : _zz_shift_i_0_10 = shift_i_map_28;
      6'b011101 : _zz_shift_i_0_10 = shift_i_map_29;
      6'b011110 : _zz_shift_i_0_10 = shift_i_map_30;
      6'b011111 : _zz_shift_i_0_10 = shift_i_map_31;
      6'b100000 : _zz_shift_i_0_10 = shift_i_map_32;
      6'b100001 : _zz_shift_i_0_10 = shift_i_map_33;
      6'b100010 : _zz_shift_i_0_10 = shift_i_map_34;
      6'b100011 : _zz_shift_i_0_10 = shift_i_map_35;
      6'b100100 : _zz_shift_i_0_10 = shift_i_map_36;
      6'b100101 : _zz_shift_i_0_10 = shift_i_map_37;
      6'b100110 : _zz_shift_i_0_10 = shift_i_map_38;
      6'b100111 : _zz_shift_i_0_10 = shift_i_map_39;
      6'b101000 : _zz_shift_i_0_10 = shift_i_map_40;
      6'b101001 : _zz_shift_i_0_10 = shift_i_map_41;
      6'b101010 : _zz_shift_i_0_10 = shift_i_map_42;
      6'b101011 : _zz_shift_i_0_10 = shift_i_map_43;
      6'b101100 : _zz_shift_i_0_10 = shift_i_map_44;
      6'b101101 : _zz_shift_i_0_10 = shift_i_map_45;
      6'b101110 : _zz_shift_i_0_10 = shift_i_map_46;
      6'b101111 : _zz_shift_i_0_10 = shift_i_map_47;
      6'b110000 : _zz_shift_i_0_10 = shift_i_map_48;
      6'b110001 : _zz_shift_i_0_10 = shift_i_map_49;
      6'b110010 : _zz_shift_i_0_10 = shift_i_map_50;
      6'b110011 : _zz_shift_i_0_10 = shift_i_map_51;
      6'b110100 : _zz_shift_i_0_10 = shift_i_map_52;
      6'b110101 : _zz_shift_i_0_10 = shift_i_map_53;
      6'b110110 : _zz_shift_i_0_10 = shift_i_map_54;
      6'b110111 : _zz_shift_i_0_10 = shift_i_map_55;
      6'b111000 : _zz_shift_i_0_10 = shift_i_map_56;
      6'b111001 : _zz_shift_i_0_10 = shift_i_map_57;
      6'b111010 : _zz_shift_i_0_10 = shift_i_map_58;
      6'b111011 : _zz_shift_i_0_10 = shift_i_map_59;
      6'b111100 : _zz_shift_i_0_10 = shift_i_map_60;
      6'b111101 : _zz_shift_i_0_10 = shift_i_map_61;
      6'b111110 : _zz_shift_i_0_10 = shift_i_map_62;
      default : _zz_shift_i_0_10 = shift_i_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_0_11)
      6'b000000 : _zz_shift_q_0_10 = shift_q_map_0;
      6'b000001 : _zz_shift_q_0_10 = shift_q_map_1;
      6'b000010 : _zz_shift_q_0_10 = shift_q_map_2;
      6'b000011 : _zz_shift_q_0_10 = shift_q_map_3;
      6'b000100 : _zz_shift_q_0_10 = shift_q_map_4;
      6'b000101 : _zz_shift_q_0_10 = shift_q_map_5;
      6'b000110 : _zz_shift_q_0_10 = shift_q_map_6;
      6'b000111 : _zz_shift_q_0_10 = shift_q_map_7;
      6'b001000 : _zz_shift_q_0_10 = shift_q_map_8;
      6'b001001 : _zz_shift_q_0_10 = shift_q_map_9;
      6'b001010 : _zz_shift_q_0_10 = shift_q_map_10;
      6'b001011 : _zz_shift_q_0_10 = shift_q_map_11;
      6'b001100 : _zz_shift_q_0_10 = shift_q_map_12;
      6'b001101 : _zz_shift_q_0_10 = shift_q_map_13;
      6'b001110 : _zz_shift_q_0_10 = shift_q_map_14;
      6'b001111 : _zz_shift_q_0_10 = shift_q_map_15;
      6'b010000 : _zz_shift_q_0_10 = shift_q_map_16;
      6'b010001 : _zz_shift_q_0_10 = shift_q_map_17;
      6'b010010 : _zz_shift_q_0_10 = shift_q_map_18;
      6'b010011 : _zz_shift_q_0_10 = shift_q_map_19;
      6'b010100 : _zz_shift_q_0_10 = shift_q_map_20;
      6'b010101 : _zz_shift_q_0_10 = shift_q_map_21;
      6'b010110 : _zz_shift_q_0_10 = shift_q_map_22;
      6'b010111 : _zz_shift_q_0_10 = shift_q_map_23;
      6'b011000 : _zz_shift_q_0_10 = shift_q_map_24;
      6'b011001 : _zz_shift_q_0_10 = shift_q_map_25;
      6'b011010 : _zz_shift_q_0_10 = shift_q_map_26;
      6'b011011 : _zz_shift_q_0_10 = shift_q_map_27;
      6'b011100 : _zz_shift_q_0_10 = shift_q_map_28;
      6'b011101 : _zz_shift_q_0_10 = shift_q_map_29;
      6'b011110 : _zz_shift_q_0_10 = shift_q_map_30;
      6'b011111 : _zz_shift_q_0_10 = shift_q_map_31;
      6'b100000 : _zz_shift_q_0_10 = shift_q_map_32;
      6'b100001 : _zz_shift_q_0_10 = shift_q_map_33;
      6'b100010 : _zz_shift_q_0_10 = shift_q_map_34;
      6'b100011 : _zz_shift_q_0_10 = shift_q_map_35;
      6'b100100 : _zz_shift_q_0_10 = shift_q_map_36;
      6'b100101 : _zz_shift_q_0_10 = shift_q_map_37;
      6'b100110 : _zz_shift_q_0_10 = shift_q_map_38;
      6'b100111 : _zz_shift_q_0_10 = shift_q_map_39;
      6'b101000 : _zz_shift_q_0_10 = shift_q_map_40;
      6'b101001 : _zz_shift_q_0_10 = shift_q_map_41;
      6'b101010 : _zz_shift_q_0_10 = shift_q_map_42;
      6'b101011 : _zz_shift_q_0_10 = shift_q_map_43;
      6'b101100 : _zz_shift_q_0_10 = shift_q_map_44;
      6'b101101 : _zz_shift_q_0_10 = shift_q_map_45;
      6'b101110 : _zz_shift_q_0_10 = shift_q_map_46;
      6'b101111 : _zz_shift_q_0_10 = shift_q_map_47;
      6'b110000 : _zz_shift_q_0_10 = shift_q_map_48;
      6'b110001 : _zz_shift_q_0_10 = shift_q_map_49;
      6'b110010 : _zz_shift_q_0_10 = shift_q_map_50;
      6'b110011 : _zz_shift_q_0_10 = shift_q_map_51;
      6'b110100 : _zz_shift_q_0_10 = shift_q_map_52;
      6'b110101 : _zz_shift_q_0_10 = shift_q_map_53;
      6'b110110 : _zz_shift_q_0_10 = shift_q_map_54;
      6'b110111 : _zz_shift_q_0_10 = shift_q_map_55;
      6'b111000 : _zz_shift_q_0_10 = shift_q_map_56;
      6'b111001 : _zz_shift_q_0_10 = shift_q_map_57;
      6'b111010 : _zz_shift_q_0_10 = shift_q_map_58;
      6'b111011 : _zz_shift_q_0_10 = shift_q_map_59;
      6'b111100 : _zz_shift_q_0_10 = shift_q_map_60;
      6'b111101 : _zz_shift_q_0_10 = shift_q_map_61;
      6'b111110 : _zz_shift_q_0_10 = shift_q_map_62;
      default : _zz_shift_q_0_10 = shift_q_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_1_11)
      6'b000000 : _zz_shift_i_1_10 = shift_i_map_0;
      6'b000001 : _zz_shift_i_1_10 = shift_i_map_1;
      6'b000010 : _zz_shift_i_1_10 = shift_i_map_2;
      6'b000011 : _zz_shift_i_1_10 = shift_i_map_3;
      6'b000100 : _zz_shift_i_1_10 = shift_i_map_4;
      6'b000101 : _zz_shift_i_1_10 = shift_i_map_5;
      6'b000110 : _zz_shift_i_1_10 = shift_i_map_6;
      6'b000111 : _zz_shift_i_1_10 = shift_i_map_7;
      6'b001000 : _zz_shift_i_1_10 = shift_i_map_8;
      6'b001001 : _zz_shift_i_1_10 = shift_i_map_9;
      6'b001010 : _zz_shift_i_1_10 = shift_i_map_10;
      6'b001011 : _zz_shift_i_1_10 = shift_i_map_11;
      6'b001100 : _zz_shift_i_1_10 = shift_i_map_12;
      6'b001101 : _zz_shift_i_1_10 = shift_i_map_13;
      6'b001110 : _zz_shift_i_1_10 = shift_i_map_14;
      6'b001111 : _zz_shift_i_1_10 = shift_i_map_15;
      6'b010000 : _zz_shift_i_1_10 = shift_i_map_16;
      6'b010001 : _zz_shift_i_1_10 = shift_i_map_17;
      6'b010010 : _zz_shift_i_1_10 = shift_i_map_18;
      6'b010011 : _zz_shift_i_1_10 = shift_i_map_19;
      6'b010100 : _zz_shift_i_1_10 = shift_i_map_20;
      6'b010101 : _zz_shift_i_1_10 = shift_i_map_21;
      6'b010110 : _zz_shift_i_1_10 = shift_i_map_22;
      6'b010111 : _zz_shift_i_1_10 = shift_i_map_23;
      6'b011000 : _zz_shift_i_1_10 = shift_i_map_24;
      6'b011001 : _zz_shift_i_1_10 = shift_i_map_25;
      6'b011010 : _zz_shift_i_1_10 = shift_i_map_26;
      6'b011011 : _zz_shift_i_1_10 = shift_i_map_27;
      6'b011100 : _zz_shift_i_1_10 = shift_i_map_28;
      6'b011101 : _zz_shift_i_1_10 = shift_i_map_29;
      6'b011110 : _zz_shift_i_1_10 = shift_i_map_30;
      6'b011111 : _zz_shift_i_1_10 = shift_i_map_31;
      6'b100000 : _zz_shift_i_1_10 = shift_i_map_32;
      6'b100001 : _zz_shift_i_1_10 = shift_i_map_33;
      6'b100010 : _zz_shift_i_1_10 = shift_i_map_34;
      6'b100011 : _zz_shift_i_1_10 = shift_i_map_35;
      6'b100100 : _zz_shift_i_1_10 = shift_i_map_36;
      6'b100101 : _zz_shift_i_1_10 = shift_i_map_37;
      6'b100110 : _zz_shift_i_1_10 = shift_i_map_38;
      6'b100111 : _zz_shift_i_1_10 = shift_i_map_39;
      6'b101000 : _zz_shift_i_1_10 = shift_i_map_40;
      6'b101001 : _zz_shift_i_1_10 = shift_i_map_41;
      6'b101010 : _zz_shift_i_1_10 = shift_i_map_42;
      6'b101011 : _zz_shift_i_1_10 = shift_i_map_43;
      6'b101100 : _zz_shift_i_1_10 = shift_i_map_44;
      6'b101101 : _zz_shift_i_1_10 = shift_i_map_45;
      6'b101110 : _zz_shift_i_1_10 = shift_i_map_46;
      6'b101111 : _zz_shift_i_1_10 = shift_i_map_47;
      6'b110000 : _zz_shift_i_1_10 = shift_i_map_48;
      6'b110001 : _zz_shift_i_1_10 = shift_i_map_49;
      6'b110010 : _zz_shift_i_1_10 = shift_i_map_50;
      6'b110011 : _zz_shift_i_1_10 = shift_i_map_51;
      6'b110100 : _zz_shift_i_1_10 = shift_i_map_52;
      6'b110101 : _zz_shift_i_1_10 = shift_i_map_53;
      6'b110110 : _zz_shift_i_1_10 = shift_i_map_54;
      6'b110111 : _zz_shift_i_1_10 = shift_i_map_55;
      6'b111000 : _zz_shift_i_1_10 = shift_i_map_56;
      6'b111001 : _zz_shift_i_1_10 = shift_i_map_57;
      6'b111010 : _zz_shift_i_1_10 = shift_i_map_58;
      6'b111011 : _zz_shift_i_1_10 = shift_i_map_59;
      6'b111100 : _zz_shift_i_1_10 = shift_i_map_60;
      6'b111101 : _zz_shift_i_1_10 = shift_i_map_61;
      6'b111110 : _zz_shift_i_1_10 = shift_i_map_62;
      default : _zz_shift_i_1_10 = shift_i_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_1_11)
      6'b000000 : _zz_shift_q_1_10 = shift_q_map_0;
      6'b000001 : _zz_shift_q_1_10 = shift_q_map_1;
      6'b000010 : _zz_shift_q_1_10 = shift_q_map_2;
      6'b000011 : _zz_shift_q_1_10 = shift_q_map_3;
      6'b000100 : _zz_shift_q_1_10 = shift_q_map_4;
      6'b000101 : _zz_shift_q_1_10 = shift_q_map_5;
      6'b000110 : _zz_shift_q_1_10 = shift_q_map_6;
      6'b000111 : _zz_shift_q_1_10 = shift_q_map_7;
      6'b001000 : _zz_shift_q_1_10 = shift_q_map_8;
      6'b001001 : _zz_shift_q_1_10 = shift_q_map_9;
      6'b001010 : _zz_shift_q_1_10 = shift_q_map_10;
      6'b001011 : _zz_shift_q_1_10 = shift_q_map_11;
      6'b001100 : _zz_shift_q_1_10 = shift_q_map_12;
      6'b001101 : _zz_shift_q_1_10 = shift_q_map_13;
      6'b001110 : _zz_shift_q_1_10 = shift_q_map_14;
      6'b001111 : _zz_shift_q_1_10 = shift_q_map_15;
      6'b010000 : _zz_shift_q_1_10 = shift_q_map_16;
      6'b010001 : _zz_shift_q_1_10 = shift_q_map_17;
      6'b010010 : _zz_shift_q_1_10 = shift_q_map_18;
      6'b010011 : _zz_shift_q_1_10 = shift_q_map_19;
      6'b010100 : _zz_shift_q_1_10 = shift_q_map_20;
      6'b010101 : _zz_shift_q_1_10 = shift_q_map_21;
      6'b010110 : _zz_shift_q_1_10 = shift_q_map_22;
      6'b010111 : _zz_shift_q_1_10 = shift_q_map_23;
      6'b011000 : _zz_shift_q_1_10 = shift_q_map_24;
      6'b011001 : _zz_shift_q_1_10 = shift_q_map_25;
      6'b011010 : _zz_shift_q_1_10 = shift_q_map_26;
      6'b011011 : _zz_shift_q_1_10 = shift_q_map_27;
      6'b011100 : _zz_shift_q_1_10 = shift_q_map_28;
      6'b011101 : _zz_shift_q_1_10 = shift_q_map_29;
      6'b011110 : _zz_shift_q_1_10 = shift_q_map_30;
      6'b011111 : _zz_shift_q_1_10 = shift_q_map_31;
      6'b100000 : _zz_shift_q_1_10 = shift_q_map_32;
      6'b100001 : _zz_shift_q_1_10 = shift_q_map_33;
      6'b100010 : _zz_shift_q_1_10 = shift_q_map_34;
      6'b100011 : _zz_shift_q_1_10 = shift_q_map_35;
      6'b100100 : _zz_shift_q_1_10 = shift_q_map_36;
      6'b100101 : _zz_shift_q_1_10 = shift_q_map_37;
      6'b100110 : _zz_shift_q_1_10 = shift_q_map_38;
      6'b100111 : _zz_shift_q_1_10 = shift_q_map_39;
      6'b101000 : _zz_shift_q_1_10 = shift_q_map_40;
      6'b101001 : _zz_shift_q_1_10 = shift_q_map_41;
      6'b101010 : _zz_shift_q_1_10 = shift_q_map_42;
      6'b101011 : _zz_shift_q_1_10 = shift_q_map_43;
      6'b101100 : _zz_shift_q_1_10 = shift_q_map_44;
      6'b101101 : _zz_shift_q_1_10 = shift_q_map_45;
      6'b101110 : _zz_shift_q_1_10 = shift_q_map_46;
      6'b101111 : _zz_shift_q_1_10 = shift_q_map_47;
      6'b110000 : _zz_shift_q_1_10 = shift_q_map_48;
      6'b110001 : _zz_shift_q_1_10 = shift_q_map_49;
      6'b110010 : _zz_shift_q_1_10 = shift_q_map_50;
      6'b110011 : _zz_shift_q_1_10 = shift_q_map_51;
      6'b110100 : _zz_shift_q_1_10 = shift_q_map_52;
      6'b110101 : _zz_shift_q_1_10 = shift_q_map_53;
      6'b110110 : _zz_shift_q_1_10 = shift_q_map_54;
      6'b110111 : _zz_shift_q_1_10 = shift_q_map_55;
      6'b111000 : _zz_shift_q_1_10 = shift_q_map_56;
      6'b111001 : _zz_shift_q_1_10 = shift_q_map_57;
      6'b111010 : _zz_shift_q_1_10 = shift_q_map_58;
      6'b111011 : _zz_shift_q_1_10 = shift_q_map_59;
      6'b111100 : _zz_shift_q_1_10 = shift_q_map_60;
      6'b111101 : _zz_shift_q_1_10 = shift_q_map_61;
      6'b111110 : _zz_shift_q_1_10 = shift_q_map_62;
      default : _zz_shift_q_1_10 = shift_q_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_2_11)
      6'b000000 : _zz_shift_i_2_10 = shift_i_map_0;
      6'b000001 : _zz_shift_i_2_10 = shift_i_map_1;
      6'b000010 : _zz_shift_i_2_10 = shift_i_map_2;
      6'b000011 : _zz_shift_i_2_10 = shift_i_map_3;
      6'b000100 : _zz_shift_i_2_10 = shift_i_map_4;
      6'b000101 : _zz_shift_i_2_10 = shift_i_map_5;
      6'b000110 : _zz_shift_i_2_10 = shift_i_map_6;
      6'b000111 : _zz_shift_i_2_10 = shift_i_map_7;
      6'b001000 : _zz_shift_i_2_10 = shift_i_map_8;
      6'b001001 : _zz_shift_i_2_10 = shift_i_map_9;
      6'b001010 : _zz_shift_i_2_10 = shift_i_map_10;
      6'b001011 : _zz_shift_i_2_10 = shift_i_map_11;
      6'b001100 : _zz_shift_i_2_10 = shift_i_map_12;
      6'b001101 : _zz_shift_i_2_10 = shift_i_map_13;
      6'b001110 : _zz_shift_i_2_10 = shift_i_map_14;
      6'b001111 : _zz_shift_i_2_10 = shift_i_map_15;
      6'b010000 : _zz_shift_i_2_10 = shift_i_map_16;
      6'b010001 : _zz_shift_i_2_10 = shift_i_map_17;
      6'b010010 : _zz_shift_i_2_10 = shift_i_map_18;
      6'b010011 : _zz_shift_i_2_10 = shift_i_map_19;
      6'b010100 : _zz_shift_i_2_10 = shift_i_map_20;
      6'b010101 : _zz_shift_i_2_10 = shift_i_map_21;
      6'b010110 : _zz_shift_i_2_10 = shift_i_map_22;
      6'b010111 : _zz_shift_i_2_10 = shift_i_map_23;
      6'b011000 : _zz_shift_i_2_10 = shift_i_map_24;
      6'b011001 : _zz_shift_i_2_10 = shift_i_map_25;
      6'b011010 : _zz_shift_i_2_10 = shift_i_map_26;
      6'b011011 : _zz_shift_i_2_10 = shift_i_map_27;
      6'b011100 : _zz_shift_i_2_10 = shift_i_map_28;
      6'b011101 : _zz_shift_i_2_10 = shift_i_map_29;
      6'b011110 : _zz_shift_i_2_10 = shift_i_map_30;
      6'b011111 : _zz_shift_i_2_10 = shift_i_map_31;
      6'b100000 : _zz_shift_i_2_10 = shift_i_map_32;
      6'b100001 : _zz_shift_i_2_10 = shift_i_map_33;
      6'b100010 : _zz_shift_i_2_10 = shift_i_map_34;
      6'b100011 : _zz_shift_i_2_10 = shift_i_map_35;
      6'b100100 : _zz_shift_i_2_10 = shift_i_map_36;
      6'b100101 : _zz_shift_i_2_10 = shift_i_map_37;
      6'b100110 : _zz_shift_i_2_10 = shift_i_map_38;
      6'b100111 : _zz_shift_i_2_10 = shift_i_map_39;
      6'b101000 : _zz_shift_i_2_10 = shift_i_map_40;
      6'b101001 : _zz_shift_i_2_10 = shift_i_map_41;
      6'b101010 : _zz_shift_i_2_10 = shift_i_map_42;
      6'b101011 : _zz_shift_i_2_10 = shift_i_map_43;
      6'b101100 : _zz_shift_i_2_10 = shift_i_map_44;
      6'b101101 : _zz_shift_i_2_10 = shift_i_map_45;
      6'b101110 : _zz_shift_i_2_10 = shift_i_map_46;
      6'b101111 : _zz_shift_i_2_10 = shift_i_map_47;
      6'b110000 : _zz_shift_i_2_10 = shift_i_map_48;
      6'b110001 : _zz_shift_i_2_10 = shift_i_map_49;
      6'b110010 : _zz_shift_i_2_10 = shift_i_map_50;
      6'b110011 : _zz_shift_i_2_10 = shift_i_map_51;
      6'b110100 : _zz_shift_i_2_10 = shift_i_map_52;
      6'b110101 : _zz_shift_i_2_10 = shift_i_map_53;
      6'b110110 : _zz_shift_i_2_10 = shift_i_map_54;
      6'b110111 : _zz_shift_i_2_10 = shift_i_map_55;
      6'b111000 : _zz_shift_i_2_10 = shift_i_map_56;
      6'b111001 : _zz_shift_i_2_10 = shift_i_map_57;
      6'b111010 : _zz_shift_i_2_10 = shift_i_map_58;
      6'b111011 : _zz_shift_i_2_10 = shift_i_map_59;
      6'b111100 : _zz_shift_i_2_10 = shift_i_map_60;
      6'b111101 : _zz_shift_i_2_10 = shift_i_map_61;
      6'b111110 : _zz_shift_i_2_10 = shift_i_map_62;
      default : _zz_shift_i_2_10 = shift_i_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_2_11)
      6'b000000 : _zz_shift_q_2_10 = shift_q_map_0;
      6'b000001 : _zz_shift_q_2_10 = shift_q_map_1;
      6'b000010 : _zz_shift_q_2_10 = shift_q_map_2;
      6'b000011 : _zz_shift_q_2_10 = shift_q_map_3;
      6'b000100 : _zz_shift_q_2_10 = shift_q_map_4;
      6'b000101 : _zz_shift_q_2_10 = shift_q_map_5;
      6'b000110 : _zz_shift_q_2_10 = shift_q_map_6;
      6'b000111 : _zz_shift_q_2_10 = shift_q_map_7;
      6'b001000 : _zz_shift_q_2_10 = shift_q_map_8;
      6'b001001 : _zz_shift_q_2_10 = shift_q_map_9;
      6'b001010 : _zz_shift_q_2_10 = shift_q_map_10;
      6'b001011 : _zz_shift_q_2_10 = shift_q_map_11;
      6'b001100 : _zz_shift_q_2_10 = shift_q_map_12;
      6'b001101 : _zz_shift_q_2_10 = shift_q_map_13;
      6'b001110 : _zz_shift_q_2_10 = shift_q_map_14;
      6'b001111 : _zz_shift_q_2_10 = shift_q_map_15;
      6'b010000 : _zz_shift_q_2_10 = shift_q_map_16;
      6'b010001 : _zz_shift_q_2_10 = shift_q_map_17;
      6'b010010 : _zz_shift_q_2_10 = shift_q_map_18;
      6'b010011 : _zz_shift_q_2_10 = shift_q_map_19;
      6'b010100 : _zz_shift_q_2_10 = shift_q_map_20;
      6'b010101 : _zz_shift_q_2_10 = shift_q_map_21;
      6'b010110 : _zz_shift_q_2_10 = shift_q_map_22;
      6'b010111 : _zz_shift_q_2_10 = shift_q_map_23;
      6'b011000 : _zz_shift_q_2_10 = shift_q_map_24;
      6'b011001 : _zz_shift_q_2_10 = shift_q_map_25;
      6'b011010 : _zz_shift_q_2_10 = shift_q_map_26;
      6'b011011 : _zz_shift_q_2_10 = shift_q_map_27;
      6'b011100 : _zz_shift_q_2_10 = shift_q_map_28;
      6'b011101 : _zz_shift_q_2_10 = shift_q_map_29;
      6'b011110 : _zz_shift_q_2_10 = shift_q_map_30;
      6'b011111 : _zz_shift_q_2_10 = shift_q_map_31;
      6'b100000 : _zz_shift_q_2_10 = shift_q_map_32;
      6'b100001 : _zz_shift_q_2_10 = shift_q_map_33;
      6'b100010 : _zz_shift_q_2_10 = shift_q_map_34;
      6'b100011 : _zz_shift_q_2_10 = shift_q_map_35;
      6'b100100 : _zz_shift_q_2_10 = shift_q_map_36;
      6'b100101 : _zz_shift_q_2_10 = shift_q_map_37;
      6'b100110 : _zz_shift_q_2_10 = shift_q_map_38;
      6'b100111 : _zz_shift_q_2_10 = shift_q_map_39;
      6'b101000 : _zz_shift_q_2_10 = shift_q_map_40;
      6'b101001 : _zz_shift_q_2_10 = shift_q_map_41;
      6'b101010 : _zz_shift_q_2_10 = shift_q_map_42;
      6'b101011 : _zz_shift_q_2_10 = shift_q_map_43;
      6'b101100 : _zz_shift_q_2_10 = shift_q_map_44;
      6'b101101 : _zz_shift_q_2_10 = shift_q_map_45;
      6'b101110 : _zz_shift_q_2_10 = shift_q_map_46;
      6'b101111 : _zz_shift_q_2_10 = shift_q_map_47;
      6'b110000 : _zz_shift_q_2_10 = shift_q_map_48;
      6'b110001 : _zz_shift_q_2_10 = shift_q_map_49;
      6'b110010 : _zz_shift_q_2_10 = shift_q_map_50;
      6'b110011 : _zz_shift_q_2_10 = shift_q_map_51;
      6'b110100 : _zz_shift_q_2_10 = shift_q_map_52;
      6'b110101 : _zz_shift_q_2_10 = shift_q_map_53;
      6'b110110 : _zz_shift_q_2_10 = shift_q_map_54;
      6'b110111 : _zz_shift_q_2_10 = shift_q_map_55;
      6'b111000 : _zz_shift_q_2_10 = shift_q_map_56;
      6'b111001 : _zz_shift_q_2_10 = shift_q_map_57;
      6'b111010 : _zz_shift_q_2_10 = shift_q_map_58;
      6'b111011 : _zz_shift_q_2_10 = shift_q_map_59;
      6'b111100 : _zz_shift_q_2_10 = shift_q_map_60;
      6'b111101 : _zz_shift_q_2_10 = shift_q_map_61;
      6'b111110 : _zz_shift_q_2_10 = shift_q_map_62;
      default : _zz_shift_q_2_10 = shift_q_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_3_11)
      6'b000000 : _zz_shift_i_3_10 = shift_i_map_0;
      6'b000001 : _zz_shift_i_3_10 = shift_i_map_1;
      6'b000010 : _zz_shift_i_3_10 = shift_i_map_2;
      6'b000011 : _zz_shift_i_3_10 = shift_i_map_3;
      6'b000100 : _zz_shift_i_3_10 = shift_i_map_4;
      6'b000101 : _zz_shift_i_3_10 = shift_i_map_5;
      6'b000110 : _zz_shift_i_3_10 = shift_i_map_6;
      6'b000111 : _zz_shift_i_3_10 = shift_i_map_7;
      6'b001000 : _zz_shift_i_3_10 = shift_i_map_8;
      6'b001001 : _zz_shift_i_3_10 = shift_i_map_9;
      6'b001010 : _zz_shift_i_3_10 = shift_i_map_10;
      6'b001011 : _zz_shift_i_3_10 = shift_i_map_11;
      6'b001100 : _zz_shift_i_3_10 = shift_i_map_12;
      6'b001101 : _zz_shift_i_3_10 = shift_i_map_13;
      6'b001110 : _zz_shift_i_3_10 = shift_i_map_14;
      6'b001111 : _zz_shift_i_3_10 = shift_i_map_15;
      6'b010000 : _zz_shift_i_3_10 = shift_i_map_16;
      6'b010001 : _zz_shift_i_3_10 = shift_i_map_17;
      6'b010010 : _zz_shift_i_3_10 = shift_i_map_18;
      6'b010011 : _zz_shift_i_3_10 = shift_i_map_19;
      6'b010100 : _zz_shift_i_3_10 = shift_i_map_20;
      6'b010101 : _zz_shift_i_3_10 = shift_i_map_21;
      6'b010110 : _zz_shift_i_3_10 = shift_i_map_22;
      6'b010111 : _zz_shift_i_3_10 = shift_i_map_23;
      6'b011000 : _zz_shift_i_3_10 = shift_i_map_24;
      6'b011001 : _zz_shift_i_3_10 = shift_i_map_25;
      6'b011010 : _zz_shift_i_3_10 = shift_i_map_26;
      6'b011011 : _zz_shift_i_3_10 = shift_i_map_27;
      6'b011100 : _zz_shift_i_3_10 = shift_i_map_28;
      6'b011101 : _zz_shift_i_3_10 = shift_i_map_29;
      6'b011110 : _zz_shift_i_3_10 = shift_i_map_30;
      6'b011111 : _zz_shift_i_3_10 = shift_i_map_31;
      6'b100000 : _zz_shift_i_3_10 = shift_i_map_32;
      6'b100001 : _zz_shift_i_3_10 = shift_i_map_33;
      6'b100010 : _zz_shift_i_3_10 = shift_i_map_34;
      6'b100011 : _zz_shift_i_3_10 = shift_i_map_35;
      6'b100100 : _zz_shift_i_3_10 = shift_i_map_36;
      6'b100101 : _zz_shift_i_3_10 = shift_i_map_37;
      6'b100110 : _zz_shift_i_3_10 = shift_i_map_38;
      6'b100111 : _zz_shift_i_3_10 = shift_i_map_39;
      6'b101000 : _zz_shift_i_3_10 = shift_i_map_40;
      6'b101001 : _zz_shift_i_3_10 = shift_i_map_41;
      6'b101010 : _zz_shift_i_3_10 = shift_i_map_42;
      6'b101011 : _zz_shift_i_3_10 = shift_i_map_43;
      6'b101100 : _zz_shift_i_3_10 = shift_i_map_44;
      6'b101101 : _zz_shift_i_3_10 = shift_i_map_45;
      6'b101110 : _zz_shift_i_3_10 = shift_i_map_46;
      6'b101111 : _zz_shift_i_3_10 = shift_i_map_47;
      6'b110000 : _zz_shift_i_3_10 = shift_i_map_48;
      6'b110001 : _zz_shift_i_3_10 = shift_i_map_49;
      6'b110010 : _zz_shift_i_3_10 = shift_i_map_50;
      6'b110011 : _zz_shift_i_3_10 = shift_i_map_51;
      6'b110100 : _zz_shift_i_3_10 = shift_i_map_52;
      6'b110101 : _zz_shift_i_3_10 = shift_i_map_53;
      6'b110110 : _zz_shift_i_3_10 = shift_i_map_54;
      6'b110111 : _zz_shift_i_3_10 = shift_i_map_55;
      6'b111000 : _zz_shift_i_3_10 = shift_i_map_56;
      6'b111001 : _zz_shift_i_3_10 = shift_i_map_57;
      6'b111010 : _zz_shift_i_3_10 = shift_i_map_58;
      6'b111011 : _zz_shift_i_3_10 = shift_i_map_59;
      6'b111100 : _zz_shift_i_3_10 = shift_i_map_60;
      6'b111101 : _zz_shift_i_3_10 = shift_i_map_61;
      6'b111110 : _zz_shift_i_3_10 = shift_i_map_62;
      default : _zz_shift_i_3_10 = shift_i_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_3_11)
      6'b000000 : _zz_shift_q_3_10 = shift_q_map_0;
      6'b000001 : _zz_shift_q_3_10 = shift_q_map_1;
      6'b000010 : _zz_shift_q_3_10 = shift_q_map_2;
      6'b000011 : _zz_shift_q_3_10 = shift_q_map_3;
      6'b000100 : _zz_shift_q_3_10 = shift_q_map_4;
      6'b000101 : _zz_shift_q_3_10 = shift_q_map_5;
      6'b000110 : _zz_shift_q_3_10 = shift_q_map_6;
      6'b000111 : _zz_shift_q_3_10 = shift_q_map_7;
      6'b001000 : _zz_shift_q_3_10 = shift_q_map_8;
      6'b001001 : _zz_shift_q_3_10 = shift_q_map_9;
      6'b001010 : _zz_shift_q_3_10 = shift_q_map_10;
      6'b001011 : _zz_shift_q_3_10 = shift_q_map_11;
      6'b001100 : _zz_shift_q_3_10 = shift_q_map_12;
      6'b001101 : _zz_shift_q_3_10 = shift_q_map_13;
      6'b001110 : _zz_shift_q_3_10 = shift_q_map_14;
      6'b001111 : _zz_shift_q_3_10 = shift_q_map_15;
      6'b010000 : _zz_shift_q_3_10 = shift_q_map_16;
      6'b010001 : _zz_shift_q_3_10 = shift_q_map_17;
      6'b010010 : _zz_shift_q_3_10 = shift_q_map_18;
      6'b010011 : _zz_shift_q_3_10 = shift_q_map_19;
      6'b010100 : _zz_shift_q_3_10 = shift_q_map_20;
      6'b010101 : _zz_shift_q_3_10 = shift_q_map_21;
      6'b010110 : _zz_shift_q_3_10 = shift_q_map_22;
      6'b010111 : _zz_shift_q_3_10 = shift_q_map_23;
      6'b011000 : _zz_shift_q_3_10 = shift_q_map_24;
      6'b011001 : _zz_shift_q_3_10 = shift_q_map_25;
      6'b011010 : _zz_shift_q_3_10 = shift_q_map_26;
      6'b011011 : _zz_shift_q_3_10 = shift_q_map_27;
      6'b011100 : _zz_shift_q_3_10 = shift_q_map_28;
      6'b011101 : _zz_shift_q_3_10 = shift_q_map_29;
      6'b011110 : _zz_shift_q_3_10 = shift_q_map_30;
      6'b011111 : _zz_shift_q_3_10 = shift_q_map_31;
      6'b100000 : _zz_shift_q_3_10 = shift_q_map_32;
      6'b100001 : _zz_shift_q_3_10 = shift_q_map_33;
      6'b100010 : _zz_shift_q_3_10 = shift_q_map_34;
      6'b100011 : _zz_shift_q_3_10 = shift_q_map_35;
      6'b100100 : _zz_shift_q_3_10 = shift_q_map_36;
      6'b100101 : _zz_shift_q_3_10 = shift_q_map_37;
      6'b100110 : _zz_shift_q_3_10 = shift_q_map_38;
      6'b100111 : _zz_shift_q_3_10 = shift_q_map_39;
      6'b101000 : _zz_shift_q_3_10 = shift_q_map_40;
      6'b101001 : _zz_shift_q_3_10 = shift_q_map_41;
      6'b101010 : _zz_shift_q_3_10 = shift_q_map_42;
      6'b101011 : _zz_shift_q_3_10 = shift_q_map_43;
      6'b101100 : _zz_shift_q_3_10 = shift_q_map_44;
      6'b101101 : _zz_shift_q_3_10 = shift_q_map_45;
      6'b101110 : _zz_shift_q_3_10 = shift_q_map_46;
      6'b101111 : _zz_shift_q_3_10 = shift_q_map_47;
      6'b110000 : _zz_shift_q_3_10 = shift_q_map_48;
      6'b110001 : _zz_shift_q_3_10 = shift_q_map_49;
      6'b110010 : _zz_shift_q_3_10 = shift_q_map_50;
      6'b110011 : _zz_shift_q_3_10 = shift_q_map_51;
      6'b110100 : _zz_shift_q_3_10 = shift_q_map_52;
      6'b110101 : _zz_shift_q_3_10 = shift_q_map_53;
      6'b110110 : _zz_shift_q_3_10 = shift_q_map_54;
      6'b110111 : _zz_shift_q_3_10 = shift_q_map_55;
      6'b111000 : _zz_shift_q_3_10 = shift_q_map_56;
      6'b111001 : _zz_shift_q_3_10 = shift_q_map_57;
      6'b111010 : _zz_shift_q_3_10 = shift_q_map_58;
      6'b111011 : _zz_shift_q_3_10 = shift_q_map_59;
      6'b111100 : _zz_shift_q_3_10 = shift_q_map_60;
      6'b111101 : _zz_shift_q_3_10 = shift_q_map_61;
      6'b111110 : _zz_shift_q_3_10 = shift_q_map_62;
      default : _zz_shift_q_3_10 = shift_q_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_4_11)
      6'b000000 : _zz_shift_i_4_10 = shift_i_map_0;
      6'b000001 : _zz_shift_i_4_10 = shift_i_map_1;
      6'b000010 : _zz_shift_i_4_10 = shift_i_map_2;
      6'b000011 : _zz_shift_i_4_10 = shift_i_map_3;
      6'b000100 : _zz_shift_i_4_10 = shift_i_map_4;
      6'b000101 : _zz_shift_i_4_10 = shift_i_map_5;
      6'b000110 : _zz_shift_i_4_10 = shift_i_map_6;
      6'b000111 : _zz_shift_i_4_10 = shift_i_map_7;
      6'b001000 : _zz_shift_i_4_10 = shift_i_map_8;
      6'b001001 : _zz_shift_i_4_10 = shift_i_map_9;
      6'b001010 : _zz_shift_i_4_10 = shift_i_map_10;
      6'b001011 : _zz_shift_i_4_10 = shift_i_map_11;
      6'b001100 : _zz_shift_i_4_10 = shift_i_map_12;
      6'b001101 : _zz_shift_i_4_10 = shift_i_map_13;
      6'b001110 : _zz_shift_i_4_10 = shift_i_map_14;
      6'b001111 : _zz_shift_i_4_10 = shift_i_map_15;
      6'b010000 : _zz_shift_i_4_10 = shift_i_map_16;
      6'b010001 : _zz_shift_i_4_10 = shift_i_map_17;
      6'b010010 : _zz_shift_i_4_10 = shift_i_map_18;
      6'b010011 : _zz_shift_i_4_10 = shift_i_map_19;
      6'b010100 : _zz_shift_i_4_10 = shift_i_map_20;
      6'b010101 : _zz_shift_i_4_10 = shift_i_map_21;
      6'b010110 : _zz_shift_i_4_10 = shift_i_map_22;
      6'b010111 : _zz_shift_i_4_10 = shift_i_map_23;
      6'b011000 : _zz_shift_i_4_10 = shift_i_map_24;
      6'b011001 : _zz_shift_i_4_10 = shift_i_map_25;
      6'b011010 : _zz_shift_i_4_10 = shift_i_map_26;
      6'b011011 : _zz_shift_i_4_10 = shift_i_map_27;
      6'b011100 : _zz_shift_i_4_10 = shift_i_map_28;
      6'b011101 : _zz_shift_i_4_10 = shift_i_map_29;
      6'b011110 : _zz_shift_i_4_10 = shift_i_map_30;
      6'b011111 : _zz_shift_i_4_10 = shift_i_map_31;
      6'b100000 : _zz_shift_i_4_10 = shift_i_map_32;
      6'b100001 : _zz_shift_i_4_10 = shift_i_map_33;
      6'b100010 : _zz_shift_i_4_10 = shift_i_map_34;
      6'b100011 : _zz_shift_i_4_10 = shift_i_map_35;
      6'b100100 : _zz_shift_i_4_10 = shift_i_map_36;
      6'b100101 : _zz_shift_i_4_10 = shift_i_map_37;
      6'b100110 : _zz_shift_i_4_10 = shift_i_map_38;
      6'b100111 : _zz_shift_i_4_10 = shift_i_map_39;
      6'b101000 : _zz_shift_i_4_10 = shift_i_map_40;
      6'b101001 : _zz_shift_i_4_10 = shift_i_map_41;
      6'b101010 : _zz_shift_i_4_10 = shift_i_map_42;
      6'b101011 : _zz_shift_i_4_10 = shift_i_map_43;
      6'b101100 : _zz_shift_i_4_10 = shift_i_map_44;
      6'b101101 : _zz_shift_i_4_10 = shift_i_map_45;
      6'b101110 : _zz_shift_i_4_10 = shift_i_map_46;
      6'b101111 : _zz_shift_i_4_10 = shift_i_map_47;
      6'b110000 : _zz_shift_i_4_10 = shift_i_map_48;
      6'b110001 : _zz_shift_i_4_10 = shift_i_map_49;
      6'b110010 : _zz_shift_i_4_10 = shift_i_map_50;
      6'b110011 : _zz_shift_i_4_10 = shift_i_map_51;
      6'b110100 : _zz_shift_i_4_10 = shift_i_map_52;
      6'b110101 : _zz_shift_i_4_10 = shift_i_map_53;
      6'b110110 : _zz_shift_i_4_10 = shift_i_map_54;
      6'b110111 : _zz_shift_i_4_10 = shift_i_map_55;
      6'b111000 : _zz_shift_i_4_10 = shift_i_map_56;
      6'b111001 : _zz_shift_i_4_10 = shift_i_map_57;
      6'b111010 : _zz_shift_i_4_10 = shift_i_map_58;
      6'b111011 : _zz_shift_i_4_10 = shift_i_map_59;
      6'b111100 : _zz_shift_i_4_10 = shift_i_map_60;
      6'b111101 : _zz_shift_i_4_10 = shift_i_map_61;
      6'b111110 : _zz_shift_i_4_10 = shift_i_map_62;
      default : _zz_shift_i_4_10 = shift_i_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_4_11)
      6'b000000 : _zz_shift_q_4_10 = shift_q_map_0;
      6'b000001 : _zz_shift_q_4_10 = shift_q_map_1;
      6'b000010 : _zz_shift_q_4_10 = shift_q_map_2;
      6'b000011 : _zz_shift_q_4_10 = shift_q_map_3;
      6'b000100 : _zz_shift_q_4_10 = shift_q_map_4;
      6'b000101 : _zz_shift_q_4_10 = shift_q_map_5;
      6'b000110 : _zz_shift_q_4_10 = shift_q_map_6;
      6'b000111 : _zz_shift_q_4_10 = shift_q_map_7;
      6'b001000 : _zz_shift_q_4_10 = shift_q_map_8;
      6'b001001 : _zz_shift_q_4_10 = shift_q_map_9;
      6'b001010 : _zz_shift_q_4_10 = shift_q_map_10;
      6'b001011 : _zz_shift_q_4_10 = shift_q_map_11;
      6'b001100 : _zz_shift_q_4_10 = shift_q_map_12;
      6'b001101 : _zz_shift_q_4_10 = shift_q_map_13;
      6'b001110 : _zz_shift_q_4_10 = shift_q_map_14;
      6'b001111 : _zz_shift_q_4_10 = shift_q_map_15;
      6'b010000 : _zz_shift_q_4_10 = shift_q_map_16;
      6'b010001 : _zz_shift_q_4_10 = shift_q_map_17;
      6'b010010 : _zz_shift_q_4_10 = shift_q_map_18;
      6'b010011 : _zz_shift_q_4_10 = shift_q_map_19;
      6'b010100 : _zz_shift_q_4_10 = shift_q_map_20;
      6'b010101 : _zz_shift_q_4_10 = shift_q_map_21;
      6'b010110 : _zz_shift_q_4_10 = shift_q_map_22;
      6'b010111 : _zz_shift_q_4_10 = shift_q_map_23;
      6'b011000 : _zz_shift_q_4_10 = shift_q_map_24;
      6'b011001 : _zz_shift_q_4_10 = shift_q_map_25;
      6'b011010 : _zz_shift_q_4_10 = shift_q_map_26;
      6'b011011 : _zz_shift_q_4_10 = shift_q_map_27;
      6'b011100 : _zz_shift_q_4_10 = shift_q_map_28;
      6'b011101 : _zz_shift_q_4_10 = shift_q_map_29;
      6'b011110 : _zz_shift_q_4_10 = shift_q_map_30;
      6'b011111 : _zz_shift_q_4_10 = shift_q_map_31;
      6'b100000 : _zz_shift_q_4_10 = shift_q_map_32;
      6'b100001 : _zz_shift_q_4_10 = shift_q_map_33;
      6'b100010 : _zz_shift_q_4_10 = shift_q_map_34;
      6'b100011 : _zz_shift_q_4_10 = shift_q_map_35;
      6'b100100 : _zz_shift_q_4_10 = shift_q_map_36;
      6'b100101 : _zz_shift_q_4_10 = shift_q_map_37;
      6'b100110 : _zz_shift_q_4_10 = shift_q_map_38;
      6'b100111 : _zz_shift_q_4_10 = shift_q_map_39;
      6'b101000 : _zz_shift_q_4_10 = shift_q_map_40;
      6'b101001 : _zz_shift_q_4_10 = shift_q_map_41;
      6'b101010 : _zz_shift_q_4_10 = shift_q_map_42;
      6'b101011 : _zz_shift_q_4_10 = shift_q_map_43;
      6'b101100 : _zz_shift_q_4_10 = shift_q_map_44;
      6'b101101 : _zz_shift_q_4_10 = shift_q_map_45;
      6'b101110 : _zz_shift_q_4_10 = shift_q_map_46;
      6'b101111 : _zz_shift_q_4_10 = shift_q_map_47;
      6'b110000 : _zz_shift_q_4_10 = shift_q_map_48;
      6'b110001 : _zz_shift_q_4_10 = shift_q_map_49;
      6'b110010 : _zz_shift_q_4_10 = shift_q_map_50;
      6'b110011 : _zz_shift_q_4_10 = shift_q_map_51;
      6'b110100 : _zz_shift_q_4_10 = shift_q_map_52;
      6'b110101 : _zz_shift_q_4_10 = shift_q_map_53;
      6'b110110 : _zz_shift_q_4_10 = shift_q_map_54;
      6'b110111 : _zz_shift_q_4_10 = shift_q_map_55;
      6'b111000 : _zz_shift_q_4_10 = shift_q_map_56;
      6'b111001 : _zz_shift_q_4_10 = shift_q_map_57;
      6'b111010 : _zz_shift_q_4_10 = shift_q_map_58;
      6'b111011 : _zz_shift_q_4_10 = shift_q_map_59;
      6'b111100 : _zz_shift_q_4_10 = shift_q_map_60;
      6'b111101 : _zz_shift_q_4_10 = shift_q_map_61;
      6'b111110 : _zz_shift_q_4_10 = shift_q_map_62;
      default : _zz_shift_q_4_10 = shift_q_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_5_11)
      6'b000000 : _zz_shift_i_5_10 = shift_i_map_0;
      6'b000001 : _zz_shift_i_5_10 = shift_i_map_1;
      6'b000010 : _zz_shift_i_5_10 = shift_i_map_2;
      6'b000011 : _zz_shift_i_5_10 = shift_i_map_3;
      6'b000100 : _zz_shift_i_5_10 = shift_i_map_4;
      6'b000101 : _zz_shift_i_5_10 = shift_i_map_5;
      6'b000110 : _zz_shift_i_5_10 = shift_i_map_6;
      6'b000111 : _zz_shift_i_5_10 = shift_i_map_7;
      6'b001000 : _zz_shift_i_5_10 = shift_i_map_8;
      6'b001001 : _zz_shift_i_5_10 = shift_i_map_9;
      6'b001010 : _zz_shift_i_5_10 = shift_i_map_10;
      6'b001011 : _zz_shift_i_5_10 = shift_i_map_11;
      6'b001100 : _zz_shift_i_5_10 = shift_i_map_12;
      6'b001101 : _zz_shift_i_5_10 = shift_i_map_13;
      6'b001110 : _zz_shift_i_5_10 = shift_i_map_14;
      6'b001111 : _zz_shift_i_5_10 = shift_i_map_15;
      6'b010000 : _zz_shift_i_5_10 = shift_i_map_16;
      6'b010001 : _zz_shift_i_5_10 = shift_i_map_17;
      6'b010010 : _zz_shift_i_5_10 = shift_i_map_18;
      6'b010011 : _zz_shift_i_5_10 = shift_i_map_19;
      6'b010100 : _zz_shift_i_5_10 = shift_i_map_20;
      6'b010101 : _zz_shift_i_5_10 = shift_i_map_21;
      6'b010110 : _zz_shift_i_5_10 = shift_i_map_22;
      6'b010111 : _zz_shift_i_5_10 = shift_i_map_23;
      6'b011000 : _zz_shift_i_5_10 = shift_i_map_24;
      6'b011001 : _zz_shift_i_5_10 = shift_i_map_25;
      6'b011010 : _zz_shift_i_5_10 = shift_i_map_26;
      6'b011011 : _zz_shift_i_5_10 = shift_i_map_27;
      6'b011100 : _zz_shift_i_5_10 = shift_i_map_28;
      6'b011101 : _zz_shift_i_5_10 = shift_i_map_29;
      6'b011110 : _zz_shift_i_5_10 = shift_i_map_30;
      6'b011111 : _zz_shift_i_5_10 = shift_i_map_31;
      6'b100000 : _zz_shift_i_5_10 = shift_i_map_32;
      6'b100001 : _zz_shift_i_5_10 = shift_i_map_33;
      6'b100010 : _zz_shift_i_5_10 = shift_i_map_34;
      6'b100011 : _zz_shift_i_5_10 = shift_i_map_35;
      6'b100100 : _zz_shift_i_5_10 = shift_i_map_36;
      6'b100101 : _zz_shift_i_5_10 = shift_i_map_37;
      6'b100110 : _zz_shift_i_5_10 = shift_i_map_38;
      6'b100111 : _zz_shift_i_5_10 = shift_i_map_39;
      6'b101000 : _zz_shift_i_5_10 = shift_i_map_40;
      6'b101001 : _zz_shift_i_5_10 = shift_i_map_41;
      6'b101010 : _zz_shift_i_5_10 = shift_i_map_42;
      6'b101011 : _zz_shift_i_5_10 = shift_i_map_43;
      6'b101100 : _zz_shift_i_5_10 = shift_i_map_44;
      6'b101101 : _zz_shift_i_5_10 = shift_i_map_45;
      6'b101110 : _zz_shift_i_5_10 = shift_i_map_46;
      6'b101111 : _zz_shift_i_5_10 = shift_i_map_47;
      6'b110000 : _zz_shift_i_5_10 = shift_i_map_48;
      6'b110001 : _zz_shift_i_5_10 = shift_i_map_49;
      6'b110010 : _zz_shift_i_5_10 = shift_i_map_50;
      6'b110011 : _zz_shift_i_5_10 = shift_i_map_51;
      6'b110100 : _zz_shift_i_5_10 = shift_i_map_52;
      6'b110101 : _zz_shift_i_5_10 = shift_i_map_53;
      6'b110110 : _zz_shift_i_5_10 = shift_i_map_54;
      6'b110111 : _zz_shift_i_5_10 = shift_i_map_55;
      6'b111000 : _zz_shift_i_5_10 = shift_i_map_56;
      6'b111001 : _zz_shift_i_5_10 = shift_i_map_57;
      6'b111010 : _zz_shift_i_5_10 = shift_i_map_58;
      6'b111011 : _zz_shift_i_5_10 = shift_i_map_59;
      6'b111100 : _zz_shift_i_5_10 = shift_i_map_60;
      6'b111101 : _zz_shift_i_5_10 = shift_i_map_61;
      6'b111110 : _zz_shift_i_5_10 = shift_i_map_62;
      default : _zz_shift_i_5_10 = shift_i_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_5_11)
      6'b000000 : _zz_shift_q_5_10 = shift_q_map_0;
      6'b000001 : _zz_shift_q_5_10 = shift_q_map_1;
      6'b000010 : _zz_shift_q_5_10 = shift_q_map_2;
      6'b000011 : _zz_shift_q_5_10 = shift_q_map_3;
      6'b000100 : _zz_shift_q_5_10 = shift_q_map_4;
      6'b000101 : _zz_shift_q_5_10 = shift_q_map_5;
      6'b000110 : _zz_shift_q_5_10 = shift_q_map_6;
      6'b000111 : _zz_shift_q_5_10 = shift_q_map_7;
      6'b001000 : _zz_shift_q_5_10 = shift_q_map_8;
      6'b001001 : _zz_shift_q_5_10 = shift_q_map_9;
      6'b001010 : _zz_shift_q_5_10 = shift_q_map_10;
      6'b001011 : _zz_shift_q_5_10 = shift_q_map_11;
      6'b001100 : _zz_shift_q_5_10 = shift_q_map_12;
      6'b001101 : _zz_shift_q_5_10 = shift_q_map_13;
      6'b001110 : _zz_shift_q_5_10 = shift_q_map_14;
      6'b001111 : _zz_shift_q_5_10 = shift_q_map_15;
      6'b010000 : _zz_shift_q_5_10 = shift_q_map_16;
      6'b010001 : _zz_shift_q_5_10 = shift_q_map_17;
      6'b010010 : _zz_shift_q_5_10 = shift_q_map_18;
      6'b010011 : _zz_shift_q_5_10 = shift_q_map_19;
      6'b010100 : _zz_shift_q_5_10 = shift_q_map_20;
      6'b010101 : _zz_shift_q_5_10 = shift_q_map_21;
      6'b010110 : _zz_shift_q_5_10 = shift_q_map_22;
      6'b010111 : _zz_shift_q_5_10 = shift_q_map_23;
      6'b011000 : _zz_shift_q_5_10 = shift_q_map_24;
      6'b011001 : _zz_shift_q_5_10 = shift_q_map_25;
      6'b011010 : _zz_shift_q_5_10 = shift_q_map_26;
      6'b011011 : _zz_shift_q_5_10 = shift_q_map_27;
      6'b011100 : _zz_shift_q_5_10 = shift_q_map_28;
      6'b011101 : _zz_shift_q_5_10 = shift_q_map_29;
      6'b011110 : _zz_shift_q_5_10 = shift_q_map_30;
      6'b011111 : _zz_shift_q_5_10 = shift_q_map_31;
      6'b100000 : _zz_shift_q_5_10 = shift_q_map_32;
      6'b100001 : _zz_shift_q_5_10 = shift_q_map_33;
      6'b100010 : _zz_shift_q_5_10 = shift_q_map_34;
      6'b100011 : _zz_shift_q_5_10 = shift_q_map_35;
      6'b100100 : _zz_shift_q_5_10 = shift_q_map_36;
      6'b100101 : _zz_shift_q_5_10 = shift_q_map_37;
      6'b100110 : _zz_shift_q_5_10 = shift_q_map_38;
      6'b100111 : _zz_shift_q_5_10 = shift_q_map_39;
      6'b101000 : _zz_shift_q_5_10 = shift_q_map_40;
      6'b101001 : _zz_shift_q_5_10 = shift_q_map_41;
      6'b101010 : _zz_shift_q_5_10 = shift_q_map_42;
      6'b101011 : _zz_shift_q_5_10 = shift_q_map_43;
      6'b101100 : _zz_shift_q_5_10 = shift_q_map_44;
      6'b101101 : _zz_shift_q_5_10 = shift_q_map_45;
      6'b101110 : _zz_shift_q_5_10 = shift_q_map_46;
      6'b101111 : _zz_shift_q_5_10 = shift_q_map_47;
      6'b110000 : _zz_shift_q_5_10 = shift_q_map_48;
      6'b110001 : _zz_shift_q_5_10 = shift_q_map_49;
      6'b110010 : _zz_shift_q_5_10 = shift_q_map_50;
      6'b110011 : _zz_shift_q_5_10 = shift_q_map_51;
      6'b110100 : _zz_shift_q_5_10 = shift_q_map_52;
      6'b110101 : _zz_shift_q_5_10 = shift_q_map_53;
      6'b110110 : _zz_shift_q_5_10 = shift_q_map_54;
      6'b110111 : _zz_shift_q_5_10 = shift_q_map_55;
      6'b111000 : _zz_shift_q_5_10 = shift_q_map_56;
      6'b111001 : _zz_shift_q_5_10 = shift_q_map_57;
      6'b111010 : _zz_shift_q_5_10 = shift_q_map_58;
      6'b111011 : _zz_shift_q_5_10 = shift_q_map_59;
      6'b111100 : _zz_shift_q_5_10 = shift_q_map_60;
      6'b111101 : _zz_shift_q_5_10 = shift_q_map_61;
      6'b111110 : _zz_shift_q_5_10 = shift_q_map_62;
      default : _zz_shift_q_5_10 = shift_q_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_6_11)
      6'b000000 : _zz_shift_i_6_10 = shift_i_map_0;
      6'b000001 : _zz_shift_i_6_10 = shift_i_map_1;
      6'b000010 : _zz_shift_i_6_10 = shift_i_map_2;
      6'b000011 : _zz_shift_i_6_10 = shift_i_map_3;
      6'b000100 : _zz_shift_i_6_10 = shift_i_map_4;
      6'b000101 : _zz_shift_i_6_10 = shift_i_map_5;
      6'b000110 : _zz_shift_i_6_10 = shift_i_map_6;
      6'b000111 : _zz_shift_i_6_10 = shift_i_map_7;
      6'b001000 : _zz_shift_i_6_10 = shift_i_map_8;
      6'b001001 : _zz_shift_i_6_10 = shift_i_map_9;
      6'b001010 : _zz_shift_i_6_10 = shift_i_map_10;
      6'b001011 : _zz_shift_i_6_10 = shift_i_map_11;
      6'b001100 : _zz_shift_i_6_10 = shift_i_map_12;
      6'b001101 : _zz_shift_i_6_10 = shift_i_map_13;
      6'b001110 : _zz_shift_i_6_10 = shift_i_map_14;
      6'b001111 : _zz_shift_i_6_10 = shift_i_map_15;
      6'b010000 : _zz_shift_i_6_10 = shift_i_map_16;
      6'b010001 : _zz_shift_i_6_10 = shift_i_map_17;
      6'b010010 : _zz_shift_i_6_10 = shift_i_map_18;
      6'b010011 : _zz_shift_i_6_10 = shift_i_map_19;
      6'b010100 : _zz_shift_i_6_10 = shift_i_map_20;
      6'b010101 : _zz_shift_i_6_10 = shift_i_map_21;
      6'b010110 : _zz_shift_i_6_10 = shift_i_map_22;
      6'b010111 : _zz_shift_i_6_10 = shift_i_map_23;
      6'b011000 : _zz_shift_i_6_10 = shift_i_map_24;
      6'b011001 : _zz_shift_i_6_10 = shift_i_map_25;
      6'b011010 : _zz_shift_i_6_10 = shift_i_map_26;
      6'b011011 : _zz_shift_i_6_10 = shift_i_map_27;
      6'b011100 : _zz_shift_i_6_10 = shift_i_map_28;
      6'b011101 : _zz_shift_i_6_10 = shift_i_map_29;
      6'b011110 : _zz_shift_i_6_10 = shift_i_map_30;
      6'b011111 : _zz_shift_i_6_10 = shift_i_map_31;
      6'b100000 : _zz_shift_i_6_10 = shift_i_map_32;
      6'b100001 : _zz_shift_i_6_10 = shift_i_map_33;
      6'b100010 : _zz_shift_i_6_10 = shift_i_map_34;
      6'b100011 : _zz_shift_i_6_10 = shift_i_map_35;
      6'b100100 : _zz_shift_i_6_10 = shift_i_map_36;
      6'b100101 : _zz_shift_i_6_10 = shift_i_map_37;
      6'b100110 : _zz_shift_i_6_10 = shift_i_map_38;
      6'b100111 : _zz_shift_i_6_10 = shift_i_map_39;
      6'b101000 : _zz_shift_i_6_10 = shift_i_map_40;
      6'b101001 : _zz_shift_i_6_10 = shift_i_map_41;
      6'b101010 : _zz_shift_i_6_10 = shift_i_map_42;
      6'b101011 : _zz_shift_i_6_10 = shift_i_map_43;
      6'b101100 : _zz_shift_i_6_10 = shift_i_map_44;
      6'b101101 : _zz_shift_i_6_10 = shift_i_map_45;
      6'b101110 : _zz_shift_i_6_10 = shift_i_map_46;
      6'b101111 : _zz_shift_i_6_10 = shift_i_map_47;
      6'b110000 : _zz_shift_i_6_10 = shift_i_map_48;
      6'b110001 : _zz_shift_i_6_10 = shift_i_map_49;
      6'b110010 : _zz_shift_i_6_10 = shift_i_map_50;
      6'b110011 : _zz_shift_i_6_10 = shift_i_map_51;
      6'b110100 : _zz_shift_i_6_10 = shift_i_map_52;
      6'b110101 : _zz_shift_i_6_10 = shift_i_map_53;
      6'b110110 : _zz_shift_i_6_10 = shift_i_map_54;
      6'b110111 : _zz_shift_i_6_10 = shift_i_map_55;
      6'b111000 : _zz_shift_i_6_10 = shift_i_map_56;
      6'b111001 : _zz_shift_i_6_10 = shift_i_map_57;
      6'b111010 : _zz_shift_i_6_10 = shift_i_map_58;
      6'b111011 : _zz_shift_i_6_10 = shift_i_map_59;
      6'b111100 : _zz_shift_i_6_10 = shift_i_map_60;
      6'b111101 : _zz_shift_i_6_10 = shift_i_map_61;
      6'b111110 : _zz_shift_i_6_10 = shift_i_map_62;
      default : _zz_shift_i_6_10 = shift_i_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_6_11)
      6'b000000 : _zz_shift_q_6_10 = shift_q_map_0;
      6'b000001 : _zz_shift_q_6_10 = shift_q_map_1;
      6'b000010 : _zz_shift_q_6_10 = shift_q_map_2;
      6'b000011 : _zz_shift_q_6_10 = shift_q_map_3;
      6'b000100 : _zz_shift_q_6_10 = shift_q_map_4;
      6'b000101 : _zz_shift_q_6_10 = shift_q_map_5;
      6'b000110 : _zz_shift_q_6_10 = shift_q_map_6;
      6'b000111 : _zz_shift_q_6_10 = shift_q_map_7;
      6'b001000 : _zz_shift_q_6_10 = shift_q_map_8;
      6'b001001 : _zz_shift_q_6_10 = shift_q_map_9;
      6'b001010 : _zz_shift_q_6_10 = shift_q_map_10;
      6'b001011 : _zz_shift_q_6_10 = shift_q_map_11;
      6'b001100 : _zz_shift_q_6_10 = shift_q_map_12;
      6'b001101 : _zz_shift_q_6_10 = shift_q_map_13;
      6'b001110 : _zz_shift_q_6_10 = shift_q_map_14;
      6'b001111 : _zz_shift_q_6_10 = shift_q_map_15;
      6'b010000 : _zz_shift_q_6_10 = shift_q_map_16;
      6'b010001 : _zz_shift_q_6_10 = shift_q_map_17;
      6'b010010 : _zz_shift_q_6_10 = shift_q_map_18;
      6'b010011 : _zz_shift_q_6_10 = shift_q_map_19;
      6'b010100 : _zz_shift_q_6_10 = shift_q_map_20;
      6'b010101 : _zz_shift_q_6_10 = shift_q_map_21;
      6'b010110 : _zz_shift_q_6_10 = shift_q_map_22;
      6'b010111 : _zz_shift_q_6_10 = shift_q_map_23;
      6'b011000 : _zz_shift_q_6_10 = shift_q_map_24;
      6'b011001 : _zz_shift_q_6_10 = shift_q_map_25;
      6'b011010 : _zz_shift_q_6_10 = shift_q_map_26;
      6'b011011 : _zz_shift_q_6_10 = shift_q_map_27;
      6'b011100 : _zz_shift_q_6_10 = shift_q_map_28;
      6'b011101 : _zz_shift_q_6_10 = shift_q_map_29;
      6'b011110 : _zz_shift_q_6_10 = shift_q_map_30;
      6'b011111 : _zz_shift_q_6_10 = shift_q_map_31;
      6'b100000 : _zz_shift_q_6_10 = shift_q_map_32;
      6'b100001 : _zz_shift_q_6_10 = shift_q_map_33;
      6'b100010 : _zz_shift_q_6_10 = shift_q_map_34;
      6'b100011 : _zz_shift_q_6_10 = shift_q_map_35;
      6'b100100 : _zz_shift_q_6_10 = shift_q_map_36;
      6'b100101 : _zz_shift_q_6_10 = shift_q_map_37;
      6'b100110 : _zz_shift_q_6_10 = shift_q_map_38;
      6'b100111 : _zz_shift_q_6_10 = shift_q_map_39;
      6'b101000 : _zz_shift_q_6_10 = shift_q_map_40;
      6'b101001 : _zz_shift_q_6_10 = shift_q_map_41;
      6'b101010 : _zz_shift_q_6_10 = shift_q_map_42;
      6'b101011 : _zz_shift_q_6_10 = shift_q_map_43;
      6'b101100 : _zz_shift_q_6_10 = shift_q_map_44;
      6'b101101 : _zz_shift_q_6_10 = shift_q_map_45;
      6'b101110 : _zz_shift_q_6_10 = shift_q_map_46;
      6'b101111 : _zz_shift_q_6_10 = shift_q_map_47;
      6'b110000 : _zz_shift_q_6_10 = shift_q_map_48;
      6'b110001 : _zz_shift_q_6_10 = shift_q_map_49;
      6'b110010 : _zz_shift_q_6_10 = shift_q_map_50;
      6'b110011 : _zz_shift_q_6_10 = shift_q_map_51;
      6'b110100 : _zz_shift_q_6_10 = shift_q_map_52;
      6'b110101 : _zz_shift_q_6_10 = shift_q_map_53;
      6'b110110 : _zz_shift_q_6_10 = shift_q_map_54;
      6'b110111 : _zz_shift_q_6_10 = shift_q_map_55;
      6'b111000 : _zz_shift_q_6_10 = shift_q_map_56;
      6'b111001 : _zz_shift_q_6_10 = shift_q_map_57;
      6'b111010 : _zz_shift_q_6_10 = shift_q_map_58;
      6'b111011 : _zz_shift_q_6_10 = shift_q_map_59;
      6'b111100 : _zz_shift_q_6_10 = shift_q_map_60;
      6'b111101 : _zz_shift_q_6_10 = shift_q_map_61;
      6'b111110 : _zz_shift_q_6_10 = shift_q_map_62;
      default : _zz_shift_q_6_10 = shift_q_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_7_11)
      6'b000000 : _zz_shift_i_7_10 = shift_i_map_0;
      6'b000001 : _zz_shift_i_7_10 = shift_i_map_1;
      6'b000010 : _zz_shift_i_7_10 = shift_i_map_2;
      6'b000011 : _zz_shift_i_7_10 = shift_i_map_3;
      6'b000100 : _zz_shift_i_7_10 = shift_i_map_4;
      6'b000101 : _zz_shift_i_7_10 = shift_i_map_5;
      6'b000110 : _zz_shift_i_7_10 = shift_i_map_6;
      6'b000111 : _zz_shift_i_7_10 = shift_i_map_7;
      6'b001000 : _zz_shift_i_7_10 = shift_i_map_8;
      6'b001001 : _zz_shift_i_7_10 = shift_i_map_9;
      6'b001010 : _zz_shift_i_7_10 = shift_i_map_10;
      6'b001011 : _zz_shift_i_7_10 = shift_i_map_11;
      6'b001100 : _zz_shift_i_7_10 = shift_i_map_12;
      6'b001101 : _zz_shift_i_7_10 = shift_i_map_13;
      6'b001110 : _zz_shift_i_7_10 = shift_i_map_14;
      6'b001111 : _zz_shift_i_7_10 = shift_i_map_15;
      6'b010000 : _zz_shift_i_7_10 = shift_i_map_16;
      6'b010001 : _zz_shift_i_7_10 = shift_i_map_17;
      6'b010010 : _zz_shift_i_7_10 = shift_i_map_18;
      6'b010011 : _zz_shift_i_7_10 = shift_i_map_19;
      6'b010100 : _zz_shift_i_7_10 = shift_i_map_20;
      6'b010101 : _zz_shift_i_7_10 = shift_i_map_21;
      6'b010110 : _zz_shift_i_7_10 = shift_i_map_22;
      6'b010111 : _zz_shift_i_7_10 = shift_i_map_23;
      6'b011000 : _zz_shift_i_7_10 = shift_i_map_24;
      6'b011001 : _zz_shift_i_7_10 = shift_i_map_25;
      6'b011010 : _zz_shift_i_7_10 = shift_i_map_26;
      6'b011011 : _zz_shift_i_7_10 = shift_i_map_27;
      6'b011100 : _zz_shift_i_7_10 = shift_i_map_28;
      6'b011101 : _zz_shift_i_7_10 = shift_i_map_29;
      6'b011110 : _zz_shift_i_7_10 = shift_i_map_30;
      6'b011111 : _zz_shift_i_7_10 = shift_i_map_31;
      6'b100000 : _zz_shift_i_7_10 = shift_i_map_32;
      6'b100001 : _zz_shift_i_7_10 = shift_i_map_33;
      6'b100010 : _zz_shift_i_7_10 = shift_i_map_34;
      6'b100011 : _zz_shift_i_7_10 = shift_i_map_35;
      6'b100100 : _zz_shift_i_7_10 = shift_i_map_36;
      6'b100101 : _zz_shift_i_7_10 = shift_i_map_37;
      6'b100110 : _zz_shift_i_7_10 = shift_i_map_38;
      6'b100111 : _zz_shift_i_7_10 = shift_i_map_39;
      6'b101000 : _zz_shift_i_7_10 = shift_i_map_40;
      6'b101001 : _zz_shift_i_7_10 = shift_i_map_41;
      6'b101010 : _zz_shift_i_7_10 = shift_i_map_42;
      6'b101011 : _zz_shift_i_7_10 = shift_i_map_43;
      6'b101100 : _zz_shift_i_7_10 = shift_i_map_44;
      6'b101101 : _zz_shift_i_7_10 = shift_i_map_45;
      6'b101110 : _zz_shift_i_7_10 = shift_i_map_46;
      6'b101111 : _zz_shift_i_7_10 = shift_i_map_47;
      6'b110000 : _zz_shift_i_7_10 = shift_i_map_48;
      6'b110001 : _zz_shift_i_7_10 = shift_i_map_49;
      6'b110010 : _zz_shift_i_7_10 = shift_i_map_50;
      6'b110011 : _zz_shift_i_7_10 = shift_i_map_51;
      6'b110100 : _zz_shift_i_7_10 = shift_i_map_52;
      6'b110101 : _zz_shift_i_7_10 = shift_i_map_53;
      6'b110110 : _zz_shift_i_7_10 = shift_i_map_54;
      6'b110111 : _zz_shift_i_7_10 = shift_i_map_55;
      6'b111000 : _zz_shift_i_7_10 = shift_i_map_56;
      6'b111001 : _zz_shift_i_7_10 = shift_i_map_57;
      6'b111010 : _zz_shift_i_7_10 = shift_i_map_58;
      6'b111011 : _zz_shift_i_7_10 = shift_i_map_59;
      6'b111100 : _zz_shift_i_7_10 = shift_i_map_60;
      6'b111101 : _zz_shift_i_7_10 = shift_i_map_61;
      6'b111110 : _zz_shift_i_7_10 = shift_i_map_62;
      default : _zz_shift_i_7_10 = shift_i_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_7_11)
      6'b000000 : _zz_shift_q_7_10 = shift_q_map_0;
      6'b000001 : _zz_shift_q_7_10 = shift_q_map_1;
      6'b000010 : _zz_shift_q_7_10 = shift_q_map_2;
      6'b000011 : _zz_shift_q_7_10 = shift_q_map_3;
      6'b000100 : _zz_shift_q_7_10 = shift_q_map_4;
      6'b000101 : _zz_shift_q_7_10 = shift_q_map_5;
      6'b000110 : _zz_shift_q_7_10 = shift_q_map_6;
      6'b000111 : _zz_shift_q_7_10 = shift_q_map_7;
      6'b001000 : _zz_shift_q_7_10 = shift_q_map_8;
      6'b001001 : _zz_shift_q_7_10 = shift_q_map_9;
      6'b001010 : _zz_shift_q_7_10 = shift_q_map_10;
      6'b001011 : _zz_shift_q_7_10 = shift_q_map_11;
      6'b001100 : _zz_shift_q_7_10 = shift_q_map_12;
      6'b001101 : _zz_shift_q_7_10 = shift_q_map_13;
      6'b001110 : _zz_shift_q_7_10 = shift_q_map_14;
      6'b001111 : _zz_shift_q_7_10 = shift_q_map_15;
      6'b010000 : _zz_shift_q_7_10 = shift_q_map_16;
      6'b010001 : _zz_shift_q_7_10 = shift_q_map_17;
      6'b010010 : _zz_shift_q_7_10 = shift_q_map_18;
      6'b010011 : _zz_shift_q_7_10 = shift_q_map_19;
      6'b010100 : _zz_shift_q_7_10 = shift_q_map_20;
      6'b010101 : _zz_shift_q_7_10 = shift_q_map_21;
      6'b010110 : _zz_shift_q_7_10 = shift_q_map_22;
      6'b010111 : _zz_shift_q_7_10 = shift_q_map_23;
      6'b011000 : _zz_shift_q_7_10 = shift_q_map_24;
      6'b011001 : _zz_shift_q_7_10 = shift_q_map_25;
      6'b011010 : _zz_shift_q_7_10 = shift_q_map_26;
      6'b011011 : _zz_shift_q_7_10 = shift_q_map_27;
      6'b011100 : _zz_shift_q_7_10 = shift_q_map_28;
      6'b011101 : _zz_shift_q_7_10 = shift_q_map_29;
      6'b011110 : _zz_shift_q_7_10 = shift_q_map_30;
      6'b011111 : _zz_shift_q_7_10 = shift_q_map_31;
      6'b100000 : _zz_shift_q_7_10 = shift_q_map_32;
      6'b100001 : _zz_shift_q_7_10 = shift_q_map_33;
      6'b100010 : _zz_shift_q_7_10 = shift_q_map_34;
      6'b100011 : _zz_shift_q_7_10 = shift_q_map_35;
      6'b100100 : _zz_shift_q_7_10 = shift_q_map_36;
      6'b100101 : _zz_shift_q_7_10 = shift_q_map_37;
      6'b100110 : _zz_shift_q_7_10 = shift_q_map_38;
      6'b100111 : _zz_shift_q_7_10 = shift_q_map_39;
      6'b101000 : _zz_shift_q_7_10 = shift_q_map_40;
      6'b101001 : _zz_shift_q_7_10 = shift_q_map_41;
      6'b101010 : _zz_shift_q_7_10 = shift_q_map_42;
      6'b101011 : _zz_shift_q_7_10 = shift_q_map_43;
      6'b101100 : _zz_shift_q_7_10 = shift_q_map_44;
      6'b101101 : _zz_shift_q_7_10 = shift_q_map_45;
      6'b101110 : _zz_shift_q_7_10 = shift_q_map_46;
      6'b101111 : _zz_shift_q_7_10 = shift_q_map_47;
      6'b110000 : _zz_shift_q_7_10 = shift_q_map_48;
      6'b110001 : _zz_shift_q_7_10 = shift_q_map_49;
      6'b110010 : _zz_shift_q_7_10 = shift_q_map_50;
      6'b110011 : _zz_shift_q_7_10 = shift_q_map_51;
      6'b110100 : _zz_shift_q_7_10 = shift_q_map_52;
      6'b110101 : _zz_shift_q_7_10 = shift_q_map_53;
      6'b110110 : _zz_shift_q_7_10 = shift_q_map_54;
      6'b110111 : _zz_shift_q_7_10 = shift_q_map_55;
      6'b111000 : _zz_shift_q_7_10 = shift_q_map_56;
      6'b111001 : _zz_shift_q_7_10 = shift_q_map_57;
      6'b111010 : _zz_shift_q_7_10 = shift_q_map_58;
      6'b111011 : _zz_shift_q_7_10 = shift_q_map_59;
      6'b111100 : _zz_shift_q_7_10 = shift_q_map_60;
      6'b111101 : _zz_shift_q_7_10 = shift_q_map_61;
      6'b111110 : _zz_shift_q_7_10 = shift_q_map_62;
      default : _zz_shift_q_7_10 = shift_q_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_0_13)
      6'b000000 : _zz_shift_i_0_12 = shift_i_map_0;
      6'b000001 : _zz_shift_i_0_12 = shift_i_map_1;
      6'b000010 : _zz_shift_i_0_12 = shift_i_map_2;
      6'b000011 : _zz_shift_i_0_12 = shift_i_map_3;
      6'b000100 : _zz_shift_i_0_12 = shift_i_map_4;
      6'b000101 : _zz_shift_i_0_12 = shift_i_map_5;
      6'b000110 : _zz_shift_i_0_12 = shift_i_map_6;
      6'b000111 : _zz_shift_i_0_12 = shift_i_map_7;
      6'b001000 : _zz_shift_i_0_12 = shift_i_map_8;
      6'b001001 : _zz_shift_i_0_12 = shift_i_map_9;
      6'b001010 : _zz_shift_i_0_12 = shift_i_map_10;
      6'b001011 : _zz_shift_i_0_12 = shift_i_map_11;
      6'b001100 : _zz_shift_i_0_12 = shift_i_map_12;
      6'b001101 : _zz_shift_i_0_12 = shift_i_map_13;
      6'b001110 : _zz_shift_i_0_12 = shift_i_map_14;
      6'b001111 : _zz_shift_i_0_12 = shift_i_map_15;
      6'b010000 : _zz_shift_i_0_12 = shift_i_map_16;
      6'b010001 : _zz_shift_i_0_12 = shift_i_map_17;
      6'b010010 : _zz_shift_i_0_12 = shift_i_map_18;
      6'b010011 : _zz_shift_i_0_12 = shift_i_map_19;
      6'b010100 : _zz_shift_i_0_12 = shift_i_map_20;
      6'b010101 : _zz_shift_i_0_12 = shift_i_map_21;
      6'b010110 : _zz_shift_i_0_12 = shift_i_map_22;
      6'b010111 : _zz_shift_i_0_12 = shift_i_map_23;
      6'b011000 : _zz_shift_i_0_12 = shift_i_map_24;
      6'b011001 : _zz_shift_i_0_12 = shift_i_map_25;
      6'b011010 : _zz_shift_i_0_12 = shift_i_map_26;
      6'b011011 : _zz_shift_i_0_12 = shift_i_map_27;
      6'b011100 : _zz_shift_i_0_12 = shift_i_map_28;
      6'b011101 : _zz_shift_i_0_12 = shift_i_map_29;
      6'b011110 : _zz_shift_i_0_12 = shift_i_map_30;
      6'b011111 : _zz_shift_i_0_12 = shift_i_map_31;
      6'b100000 : _zz_shift_i_0_12 = shift_i_map_32;
      6'b100001 : _zz_shift_i_0_12 = shift_i_map_33;
      6'b100010 : _zz_shift_i_0_12 = shift_i_map_34;
      6'b100011 : _zz_shift_i_0_12 = shift_i_map_35;
      6'b100100 : _zz_shift_i_0_12 = shift_i_map_36;
      6'b100101 : _zz_shift_i_0_12 = shift_i_map_37;
      6'b100110 : _zz_shift_i_0_12 = shift_i_map_38;
      6'b100111 : _zz_shift_i_0_12 = shift_i_map_39;
      6'b101000 : _zz_shift_i_0_12 = shift_i_map_40;
      6'b101001 : _zz_shift_i_0_12 = shift_i_map_41;
      6'b101010 : _zz_shift_i_0_12 = shift_i_map_42;
      6'b101011 : _zz_shift_i_0_12 = shift_i_map_43;
      6'b101100 : _zz_shift_i_0_12 = shift_i_map_44;
      6'b101101 : _zz_shift_i_0_12 = shift_i_map_45;
      6'b101110 : _zz_shift_i_0_12 = shift_i_map_46;
      6'b101111 : _zz_shift_i_0_12 = shift_i_map_47;
      6'b110000 : _zz_shift_i_0_12 = shift_i_map_48;
      6'b110001 : _zz_shift_i_0_12 = shift_i_map_49;
      6'b110010 : _zz_shift_i_0_12 = shift_i_map_50;
      6'b110011 : _zz_shift_i_0_12 = shift_i_map_51;
      6'b110100 : _zz_shift_i_0_12 = shift_i_map_52;
      6'b110101 : _zz_shift_i_0_12 = shift_i_map_53;
      6'b110110 : _zz_shift_i_0_12 = shift_i_map_54;
      6'b110111 : _zz_shift_i_0_12 = shift_i_map_55;
      6'b111000 : _zz_shift_i_0_12 = shift_i_map_56;
      6'b111001 : _zz_shift_i_0_12 = shift_i_map_57;
      6'b111010 : _zz_shift_i_0_12 = shift_i_map_58;
      6'b111011 : _zz_shift_i_0_12 = shift_i_map_59;
      6'b111100 : _zz_shift_i_0_12 = shift_i_map_60;
      6'b111101 : _zz_shift_i_0_12 = shift_i_map_61;
      6'b111110 : _zz_shift_i_0_12 = shift_i_map_62;
      default : _zz_shift_i_0_12 = shift_i_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_0_13)
      6'b000000 : _zz_shift_q_0_12 = shift_q_map_0;
      6'b000001 : _zz_shift_q_0_12 = shift_q_map_1;
      6'b000010 : _zz_shift_q_0_12 = shift_q_map_2;
      6'b000011 : _zz_shift_q_0_12 = shift_q_map_3;
      6'b000100 : _zz_shift_q_0_12 = shift_q_map_4;
      6'b000101 : _zz_shift_q_0_12 = shift_q_map_5;
      6'b000110 : _zz_shift_q_0_12 = shift_q_map_6;
      6'b000111 : _zz_shift_q_0_12 = shift_q_map_7;
      6'b001000 : _zz_shift_q_0_12 = shift_q_map_8;
      6'b001001 : _zz_shift_q_0_12 = shift_q_map_9;
      6'b001010 : _zz_shift_q_0_12 = shift_q_map_10;
      6'b001011 : _zz_shift_q_0_12 = shift_q_map_11;
      6'b001100 : _zz_shift_q_0_12 = shift_q_map_12;
      6'b001101 : _zz_shift_q_0_12 = shift_q_map_13;
      6'b001110 : _zz_shift_q_0_12 = shift_q_map_14;
      6'b001111 : _zz_shift_q_0_12 = shift_q_map_15;
      6'b010000 : _zz_shift_q_0_12 = shift_q_map_16;
      6'b010001 : _zz_shift_q_0_12 = shift_q_map_17;
      6'b010010 : _zz_shift_q_0_12 = shift_q_map_18;
      6'b010011 : _zz_shift_q_0_12 = shift_q_map_19;
      6'b010100 : _zz_shift_q_0_12 = shift_q_map_20;
      6'b010101 : _zz_shift_q_0_12 = shift_q_map_21;
      6'b010110 : _zz_shift_q_0_12 = shift_q_map_22;
      6'b010111 : _zz_shift_q_0_12 = shift_q_map_23;
      6'b011000 : _zz_shift_q_0_12 = shift_q_map_24;
      6'b011001 : _zz_shift_q_0_12 = shift_q_map_25;
      6'b011010 : _zz_shift_q_0_12 = shift_q_map_26;
      6'b011011 : _zz_shift_q_0_12 = shift_q_map_27;
      6'b011100 : _zz_shift_q_0_12 = shift_q_map_28;
      6'b011101 : _zz_shift_q_0_12 = shift_q_map_29;
      6'b011110 : _zz_shift_q_0_12 = shift_q_map_30;
      6'b011111 : _zz_shift_q_0_12 = shift_q_map_31;
      6'b100000 : _zz_shift_q_0_12 = shift_q_map_32;
      6'b100001 : _zz_shift_q_0_12 = shift_q_map_33;
      6'b100010 : _zz_shift_q_0_12 = shift_q_map_34;
      6'b100011 : _zz_shift_q_0_12 = shift_q_map_35;
      6'b100100 : _zz_shift_q_0_12 = shift_q_map_36;
      6'b100101 : _zz_shift_q_0_12 = shift_q_map_37;
      6'b100110 : _zz_shift_q_0_12 = shift_q_map_38;
      6'b100111 : _zz_shift_q_0_12 = shift_q_map_39;
      6'b101000 : _zz_shift_q_0_12 = shift_q_map_40;
      6'b101001 : _zz_shift_q_0_12 = shift_q_map_41;
      6'b101010 : _zz_shift_q_0_12 = shift_q_map_42;
      6'b101011 : _zz_shift_q_0_12 = shift_q_map_43;
      6'b101100 : _zz_shift_q_0_12 = shift_q_map_44;
      6'b101101 : _zz_shift_q_0_12 = shift_q_map_45;
      6'b101110 : _zz_shift_q_0_12 = shift_q_map_46;
      6'b101111 : _zz_shift_q_0_12 = shift_q_map_47;
      6'b110000 : _zz_shift_q_0_12 = shift_q_map_48;
      6'b110001 : _zz_shift_q_0_12 = shift_q_map_49;
      6'b110010 : _zz_shift_q_0_12 = shift_q_map_50;
      6'b110011 : _zz_shift_q_0_12 = shift_q_map_51;
      6'b110100 : _zz_shift_q_0_12 = shift_q_map_52;
      6'b110101 : _zz_shift_q_0_12 = shift_q_map_53;
      6'b110110 : _zz_shift_q_0_12 = shift_q_map_54;
      6'b110111 : _zz_shift_q_0_12 = shift_q_map_55;
      6'b111000 : _zz_shift_q_0_12 = shift_q_map_56;
      6'b111001 : _zz_shift_q_0_12 = shift_q_map_57;
      6'b111010 : _zz_shift_q_0_12 = shift_q_map_58;
      6'b111011 : _zz_shift_q_0_12 = shift_q_map_59;
      6'b111100 : _zz_shift_q_0_12 = shift_q_map_60;
      6'b111101 : _zz_shift_q_0_12 = shift_q_map_61;
      6'b111110 : _zz_shift_q_0_12 = shift_q_map_62;
      default : _zz_shift_q_0_12 = shift_q_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_1_13)
      6'b000000 : _zz_shift_i_1_12 = shift_i_map_0;
      6'b000001 : _zz_shift_i_1_12 = shift_i_map_1;
      6'b000010 : _zz_shift_i_1_12 = shift_i_map_2;
      6'b000011 : _zz_shift_i_1_12 = shift_i_map_3;
      6'b000100 : _zz_shift_i_1_12 = shift_i_map_4;
      6'b000101 : _zz_shift_i_1_12 = shift_i_map_5;
      6'b000110 : _zz_shift_i_1_12 = shift_i_map_6;
      6'b000111 : _zz_shift_i_1_12 = shift_i_map_7;
      6'b001000 : _zz_shift_i_1_12 = shift_i_map_8;
      6'b001001 : _zz_shift_i_1_12 = shift_i_map_9;
      6'b001010 : _zz_shift_i_1_12 = shift_i_map_10;
      6'b001011 : _zz_shift_i_1_12 = shift_i_map_11;
      6'b001100 : _zz_shift_i_1_12 = shift_i_map_12;
      6'b001101 : _zz_shift_i_1_12 = shift_i_map_13;
      6'b001110 : _zz_shift_i_1_12 = shift_i_map_14;
      6'b001111 : _zz_shift_i_1_12 = shift_i_map_15;
      6'b010000 : _zz_shift_i_1_12 = shift_i_map_16;
      6'b010001 : _zz_shift_i_1_12 = shift_i_map_17;
      6'b010010 : _zz_shift_i_1_12 = shift_i_map_18;
      6'b010011 : _zz_shift_i_1_12 = shift_i_map_19;
      6'b010100 : _zz_shift_i_1_12 = shift_i_map_20;
      6'b010101 : _zz_shift_i_1_12 = shift_i_map_21;
      6'b010110 : _zz_shift_i_1_12 = shift_i_map_22;
      6'b010111 : _zz_shift_i_1_12 = shift_i_map_23;
      6'b011000 : _zz_shift_i_1_12 = shift_i_map_24;
      6'b011001 : _zz_shift_i_1_12 = shift_i_map_25;
      6'b011010 : _zz_shift_i_1_12 = shift_i_map_26;
      6'b011011 : _zz_shift_i_1_12 = shift_i_map_27;
      6'b011100 : _zz_shift_i_1_12 = shift_i_map_28;
      6'b011101 : _zz_shift_i_1_12 = shift_i_map_29;
      6'b011110 : _zz_shift_i_1_12 = shift_i_map_30;
      6'b011111 : _zz_shift_i_1_12 = shift_i_map_31;
      6'b100000 : _zz_shift_i_1_12 = shift_i_map_32;
      6'b100001 : _zz_shift_i_1_12 = shift_i_map_33;
      6'b100010 : _zz_shift_i_1_12 = shift_i_map_34;
      6'b100011 : _zz_shift_i_1_12 = shift_i_map_35;
      6'b100100 : _zz_shift_i_1_12 = shift_i_map_36;
      6'b100101 : _zz_shift_i_1_12 = shift_i_map_37;
      6'b100110 : _zz_shift_i_1_12 = shift_i_map_38;
      6'b100111 : _zz_shift_i_1_12 = shift_i_map_39;
      6'b101000 : _zz_shift_i_1_12 = shift_i_map_40;
      6'b101001 : _zz_shift_i_1_12 = shift_i_map_41;
      6'b101010 : _zz_shift_i_1_12 = shift_i_map_42;
      6'b101011 : _zz_shift_i_1_12 = shift_i_map_43;
      6'b101100 : _zz_shift_i_1_12 = shift_i_map_44;
      6'b101101 : _zz_shift_i_1_12 = shift_i_map_45;
      6'b101110 : _zz_shift_i_1_12 = shift_i_map_46;
      6'b101111 : _zz_shift_i_1_12 = shift_i_map_47;
      6'b110000 : _zz_shift_i_1_12 = shift_i_map_48;
      6'b110001 : _zz_shift_i_1_12 = shift_i_map_49;
      6'b110010 : _zz_shift_i_1_12 = shift_i_map_50;
      6'b110011 : _zz_shift_i_1_12 = shift_i_map_51;
      6'b110100 : _zz_shift_i_1_12 = shift_i_map_52;
      6'b110101 : _zz_shift_i_1_12 = shift_i_map_53;
      6'b110110 : _zz_shift_i_1_12 = shift_i_map_54;
      6'b110111 : _zz_shift_i_1_12 = shift_i_map_55;
      6'b111000 : _zz_shift_i_1_12 = shift_i_map_56;
      6'b111001 : _zz_shift_i_1_12 = shift_i_map_57;
      6'b111010 : _zz_shift_i_1_12 = shift_i_map_58;
      6'b111011 : _zz_shift_i_1_12 = shift_i_map_59;
      6'b111100 : _zz_shift_i_1_12 = shift_i_map_60;
      6'b111101 : _zz_shift_i_1_12 = shift_i_map_61;
      6'b111110 : _zz_shift_i_1_12 = shift_i_map_62;
      default : _zz_shift_i_1_12 = shift_i_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_1_13)
      6'b000000 : _zz_shift_q_1_12 = shift_q_map_0;
      6'b000001 : _zz_shift_q_1_12 = shift_q_map_1;
      6'b000010 : _zz_shift_q_1_12 = shift_q_map_2;
      6'b000011 : _zz_shift_q_1_12 = shift_q_map_3;
      6'b000100 : _zz_shift_q_1_12 = shift_q_map_4;
      6'b000101 : _zz_shift_q_1_12 = shift_q_map_5;
      6'b000110 : _zz_shift_q_1_12 = shift_q_map_6;
      6'b000111 : _zz_shift_q_1_12 = shift_q_map_7;
      6'b001000 : _zz_shift_q_1_12 = shift_q_map_8;
      6'b001001 : _zz_shift_q_1_12 = shift_q_map_9;
      6'b001010 : _zz_shift_q_1_12 = shift_q_map_10;
      6'b001011 : _zz_shift_q_1_12 = shift_q_map_11;
      6'b001100 : _zz_shift_q_1_12 = shift_q_map_12;
      6'b001101 : _zz_shift_q_1_12 = shift_q_map_13;
      6'b001110 : _zz_shift_q_1_12 = shift_q_map_14;
      6'b001111 : _zz_shift_q_1_12 = shift_q_map_15;
      6'b010000 : _zz_shift_q_1_12 = shift_q_map_16;
      6'b010001 : _zz_shift_q_1_12 = shift_q_map_17;
      6'b010010 : _zz_shift_q_1_12 = shift_q_map_18;
      6'b010011 : _zz_shift_q_1_12 = shift_q_map_19;
      6'b010100 : _zz_shift_q_1_12 = shift_q_map_20;
      6'b010101 : _zz_shift_q_1_12 = shift_q_map_21;
      6'b010110 : _zz_shift_q_1_12 = shift_q_map_22;
      6'b010111 : _zz_shift_q_1_12 = shift_q_map_23;
      6'b011000 : _zz_shift_q_1_12 = shift_q_map_24;
      6'b011001 : _zz_shift_q_1_12 = shift_q_map_25;
      6'b011010 : _zz_shift_q_1_12 = shift_q_map_26;
      6'b011011 : _zz_shift_q_1_12 = shift_q_map_27;
      6'b011100 : _zz_shift_q_1_12 = shift_q_map_28;
      6'b011101 : _zz_shift_q_1_12 = shift_q_map_29;
      6'b011110 : _zz_shift_q_1_12 = shift_q_map_30;
      6'b011111 : _zz_shift_q_1_12 = shift_q_map_31;
      6'b100000 : _zz_shift_q_1_12 = shift_q_map_32;
      6'b100001 : _zz_shift_q_1_12 = shift_q_map_33;
      6'b100010 : _zz_shift_q_1_12 = shift_q_map_34;
      6'b100011 : _zz_shift_q_1_12 = shift_q_map_35;
      6'b100100 : _zz_shift_q_1_12 = shift_q_map_36;
      6'b100101 : _zz_shift_q_1_12 = shift_q_map_37;
      6'b100110 : _zz_shift_q_1_12 = shift_q_map_38;
      6'b100111 : _zz_shift_q_1_12 = shift_q_map_39;
      6'b101000 : _zz_shift_q_1_12 = shift_q_map_40;
      6'b101001 : _zz_shift_q_1_12 = shift_q_map_41;
      6'b101010 : _zz_shift_q_1_12 = shift_q_map_42;
      6'b101011 : _zz_shift_q_1_12 = shift_q_map_43;
      6'b101100 : _zz_shift_q_1_12 = shift_q_map_44;
      6'b101101 : _zz_shift_q_1_12 = shift_q_map_45;
      6'b101110 : _zz_shift_q_1_12 = shift_q_map_46;
      6'b101111 : _zz_shift_q_1_12 = shift_q_map_47;
      6'b110000 : _zz_shift_q_1_12 = shift_q_map_48;
      6'b110001 : _zz_shift_q_1_12 = shift_q_map_49;
      6'b110010 : _zz_shift_q_1_12 = shift_q_map_50;
      6'b110011 : _zz_shift_q_1_12 = shift_q_map_51;
      6'b110100 : _zz_shift_q_1_12 = shift_q_map_52;
      6'b110101 : _zz_shift_q_1_12 = shift_q_map_53;
      6'b110110 : _zz_shift_q_1_12 = shift_q_map_54;
      6'b110111 : _zz_shift_q_1_12 = shift_q_map_55;
      6'b111000 : _zz_shift_q_1_12 = shift_q_map_56;
      6'b111001 : _zz_shift_q_1_12 = shift_q_map_57;
      6'b111010 : _zz_shift_q_1_12 = shift_q_map_58;
      6'b111011 : _zz_shift_q_1_12 = shift_q_map_59;
      6'b111100 : _zz_shift_q_1_12 = shift_q_map_60;
      6'b111101 : _zz_shift_q_1_12 = shift_q_map_61;
      6'b111110 : _zz_shift_q_1_12 = shift_q_map_62;
      default : _zz_shift_q_1_12 = shift_q_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_2_13)
      6'b000000 : _zz_shift_i_2_12 = shift_i_map_0;
      6'b000001 : _zz_shift_i_2_12 = shift_i_map_1;
      6'b000010 : _zz_shift_i_2_12 = shift_i_map_2;
      6'b000011 : _zz_shift_i_2_12 = shift_i_map_3;
      6'b000100 : _zz_shift_i_2_12 = shift_i_map_4;
      6'b000101 : _zz_shift_i_2_12 = shift_i_map_5;
      6'b000110 : _zz_shift_i_2_12 = shift_i_map_6;
      6'b000111 : _zz_shift_i_2_12 = shift_i_map_7;
      6'b001000 : _zz_shift_i_2_12 = shift_i_map_8;
      6'b001001 : _zz_shift_i_2_12 = shift_i_map_9;
      6'b001010 : _zz_shift_i_2_12 = shift_i_map_10;
      6'b001011 : _zz_shift_i_2_12 = shift_i_map_11;
      6'b001100 : _zz_shift_i_2_12 = shift_i_map_12;
      6'b001101 : _zz_shift_i_2_12 = shift_i_map_13;
      6'b001110 : _zz_shift_i_2_12 = shift_i_map_14;
      6'b001111 : _zz_shift_i_2_12 = shift_i_map_15;
      6'b010000 : _zz_shift_i_2_12 = shift_i_map_16;
      6'b010001 : _zz_shift_i_2_12 = shift_i_map_17;
      6'b010010 : _zz_shift_i_2_12 = shift_i_map_18;
      6'b010011 : _zz_shift_i_2_12 = shift_i_map_19;
      6'b010100 : _zz_shift_i_2_12 = shift_i_map_20;
      6'b010101 : _zz_shift_i_2_12 = shift_i_map_21;
      6'b010110 : _zz_shift_i_2_12 = shift_i_map_22;
      6'b010111 : _zz_shift_i_2_12 = shift_i_map_23;
      6'b011000 : _zz_shift_i_2_12 = shift_i_map_24;
      6'b011001 : _zz_shift_i_2_12 = shift_i_map_25;
      6'b011010 : _zz_shift_i_2_12 = shift_i_map_26;
      6'b011011 : _zz_shift_i_2_12 = shift_i_map_27;
      6'b011100 : _zz_shift_i_2_12 = shift_i_map_28;
      6'b011101 : _zz_shift_i_2_12 = shift_i_map_29;
      6'b011110 : _zz_shift_i_2_12 = shift_i_map_30;
      6'b011111 : _zz_shift_i_2_12 = shift_i_map_31;
      6'b100000 : _zz_shift_i_2_12 = shift_i_map_32;
      6'b100001 : _zz_shift_i_2_12 = shift_i_map_33;
      6'b100010 : _zz_shift_i_2_12 = shift_i_map_34;
      6'b100011 : _zz_shift_i_2_12 = shift_i_map_35;
      6'b100100 : _zz_shift_i_2_12 = shift_i_map_36;
      6'b100101 : _zz_shift_i_2_12 = shift_i_map_37;
      6'b100110 : _zz_shift_i_2_12 = shift_i_map_38;
      6'b100111 : _zz_shift_i_2_12 = shift_i_map_39;
      6'b101000 : _zz_shift_i_2_12 = shift_i_map_40;
      6'b101001 : _zz_shift_i_2_12 = shift_i_map_41;
      6'b101010 : _zz_shift_i_2_12 = shift_i_map_42;
      6'b101011 : _zz_shift_i_2_12 = shift_i_map_43;
      6'b101100 : _zz_shift_i_2_12 = shift_i_map_44;
      6'b101101 : _zz_shift_i_2_12 = shift_i_map_45;
      6'b101110 : _zz_shift_i_2_12 = shift_i_map_46;
      6'b101111 : _zz_shift_i_2_12 = shift_i_map_47;
      6'b110000 : _zz_shift_i_2_12 = shift_i_map_48;
      6'b110001 : _zz_shift_i_2_12 = shift_i_map_49;
      6'b110010 : _zz_shift_i_2_12 = shift_i_map_50;
      6'b110011 : _zz_shift_i_2_12 = shift_i_map_51;
      6'b110100 : _zz_shift_i_2_12 = shift_i_map_52;
      6'b110101 : _zz_shift_i_2_12 = shift_i_map_53;
      6'b110110 : _zz_shift_i_2_12 = shift_i_map_54;
      6'b110111 : _zz_shift_i_2_12 = shift_i_map_55;
      6'b111000 : _zz_shift_i_2_12 = shift_i_map_56;
      6'b111001 : _zz_shift_i_2_12 = shift_i_map_57;
      6'b111010 : _zz_shift_i_2_12 = shift_i_map_58;
      6'b111011 : _zz_shift_i_2_12 = shift_i_map_59;
      6'b111100 : _zz_shift_i_2_12 = shift_i_map_60;
      6'b111101 : _zz_shift_i_2_12 = shift_i_map_61;
      6'b111110 : _zz_shift_i_2_12 = shift_i_map_62;
      default : _zz_shift_i_2_12 = shift_i_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_2_13)
      6'b000000 : _zz_shift_q_2_12 = shift_q_map_0;
      6'b000001 : _zz_shift_q_2_12 = shift_q_map_1;
      6'b000010 : _zz_shift_q_2_12 = shift_q_map_2;
      6'b000011 : _zz_shift_q_2_12 = shift_q_map_3;
      6'b000100 : _zz_shift_q_2_12 = shift_q_map_4;
      6'b000101 : _zz_shift_q_2_12 = shift_q_map_5;
      6'b000110 : _zz_shift_q_2_12 = shift_q_map_6;
      6'b000111 : _zz_shift_q_2_12 = shift_q_map_7;
      6'b001000 : _zz_shift_q_2_12 = shift_q_map_8;
      6'b001001 : _zz_shift_q_2_12 = shift_q_map_9;
      6'b001010 : _zz_shift_q_2_12 = shift_q_map_10;
      6'b001011 : _zz_shift_q_2_12 = shift_q_map_11;
      6'b001100 : _zz_shift_q_2_12 = shift_q_map_12;
      6'b001101 : _zz_shift_q_2_12 = shift_q_map_13;
      6'b001110 : _zz_shift_q_2_12 = shift_q_map_14;
      6'b001111 : _zz_shift_q_2_12 = shift_q_map_15;
      6'b010000 : _zz_shift_q_2_12 = shift_q_map_16;
      6'b010001 : _zz_shift_q_2_12 = shift_q_map_17;
      6'b010010 : _zz_shift_q_2_12 = shift_q_map_18;
      6'b010011 : _zz_shift_q_2_12 = shift_q_map_19;
      6'b010100 : _zz_shift_q_2_12 = shift_q_map_20;
      6'b010101 : _zz_shift_q_2_12 = shift_q_map_21;
      6'b010110 : _zz_shift_q_2_12 = shift_q_map_22;
      6'b010111 : _zz_shift_q_2_12 = shift_q_map_23;
      6'b011000 : _zz_shift_q_2_12 = shift_q_map_24;
      6'b011001 : _zz_shift_q_2_12 = shift_q_map_25;
      6'b011010 : _zz_shift_q_2_12 = shift_q_map_26;
      6'b011011 : _zz_shift_q_2_12 = shift_q_map_27;
      6'b011100 : _zz_shift_q_2_12 = shift_q_map_28;
      6'b011101 : _zz_shift_q_2_12 = shift_q_map_29;
      6'b011110 : _zz_shift_q_2_12 = shift_q_map_30;
      6'b011111 : _zz_shift_q_2_12 = shift_q_map_31;
      6'b100000 : _zz_shift_q_2_12 = shift_q_map_32;
      6'b100001 : _zz_shift_q_2_12 = shift_q_map_33;
      6'b100010 : _zz_shift_q_2_12 = shift_q_map_34;
      6'b100011 : _zz_shift_q_2_12 = shift_q_map_35;
      6'b100100 : _zz_shift_q_2_12 = shift_q_map_36;
      6'b100101 : _zz_shift_q_2_12 = shift_q_map_37;
      6'b100110 : _zz_shift_q_2_12 = shift_q_map_38;
      6'b100111 : _zz_shift_q_2_12 = shift_q_map_39;
      6'b101000 : _zz_shift_q_2_12 = shift_q_map_40;
      6'b101001 : _zz_shift_q_2_12 = shift_q_map_41;
      6'b101010 : _zz_shift_q_2_12 = shift_q_map_42;
      6'b101011 : _zz_shift_q_2_12 = shift_q_map_43;
      6'b101100 : _zz_shift_q_2_12 = shift_q_map_44;
      6'b101101 : _zz_shift_q_2_12 = shift_q_map_45;
      6'b101110 : _zz_shift_q_2_12 = shift_q_map_46;
      6'b101111 : _zz_shift_q_2_12 = shift_q_map_47;
      6'b110000 : _zz_shift_q_2_12 = shift_q_map_48;
      6'b110001 : _zz_shift_q_2_12 = shift_q_map_49;
      6'b110010 : _zz_shift_q_2_12 = shift_q_map_50;
      6'b110011 : _zz_shift_q_2_12 = shift_q_map_51;
      6'b110100 : _zz_shift_q_2_12 = shift_q_map_52;
      6'b110101 : _zz_shift_q_2_12 = shift_q_map_53;
      6'b110110 : _zz_shift_q_2_12 = shift_q_map_54;
      6'b110111 : _zz_shift_q_2_12 = shift_q_map_55;
      6'b111000 : _zz_shift_q_2_12 = shift_q_map_56;
      6'b111001 : _zz_shift_q_2_12 = shift_q_map_57;
      6'b111010 : _zz_shift_q_2_12 = shift_q_map_58;
      6'b111011 : _zz_shift_q_2_12 = shift_q_map_59;
      6'b111100 : _zz_shift_q_2_12 = shift_q_map_60;
      6'b111101 : _zz_shift_q_2_12 = shift_q_map_61;
      6'b111110 : _zz_shift_q_2_12 = shift_q_map_62;
      default : _zz_shift_q_2_12 = shift_q_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_3_13)
      6'b000000 : _zz_shift_i_3_12 = shift_i_map_0;
      6'b000001 : _zz_shift_i_3_12 = shift_i_map_1;
      6'b000010 : _zz_shift_i_3_12 = shift_i_map_2;
      6'b000011 : _zz_shift_i_3_12 = shift_i_map_3;
      6'b000100 : _zz_shift_i_3_12 = shift_i_map_4;
      6'b000101 : _zz_shift_i_3_12 = shift_i_map_5;
      6'b000110 : _zz_shift_i_3_12 = shift_i_map_6;
      6'b000111 : _zz_shift_i_3_12 = shift_i_map_7;
      6'b001000 : _zz_shift_i_3_12 = shift_i_map_8;
      6'b001001 : _zz_shift_i_3_12 = shift_i_map_9;
      6'b001010 : _zz_shift_i_3_12 = shift_i_map_10;
      6'b001011 : _zz_shift_i_3_12 = shift_i_map_11;
      6'b001100 : _zz_shift_i_3_12 = shift_i_map_12;
      6'b001101 : _zz_shift_i_3_12 = shift_i_map_13;
      6'b001110 : _zz_shift_i_3_12 = shift_i_map_14;
      6'b001111 : _zz_shift_i_3_12 = shift_i_map_15;
      6'b010000 : _zz_shift_i_3_12 = shift_i_map_16;
      6'b010001 : _zz_shift_i_3_12 = shift_i_map_17;
      6'b010010 : _zz_shift_i_3_12 = shift_i_map_18;
      6'b010011 : _zz_shift_i_3_12 = shift_i_map_19;
      6'b010100 : _zz_shift_i_3_12 = shift_i_map_20;
      6'b010101 : _zz_shift_i_3_12 = shift_i_map_21;
      6'b010110 : _zz_shift_i_3_12 = shift_i_map_22;
      6'b010111 : _zz_shift_i_3_12 = shift_i_map_23;
      6'b011000 : _zz_shift_i_3_12 = shift_i_map_24;
      6'b011001 : _zz_shift_i_3_12 = shift_i_map_25;
      6'b011010 : _zz_shift_i_3_12 = shift_i_map_26;
      6'b011011 : _zz_shift_i_3_12 = shift_i_map_27;
      6'b011100 : _zz_shift_i_3_12 = shift_i_map_28;
      6'b011101 : _zz_shift_i_3_12 = shift_i_map_29;
      6'b011110 : _zz_shift_i_3_12 = shift_i_map_30;
      6'b011111 : _zz_shift_i_3_12 = shift_i_map_31;
      6'b100000 : _zz_shift_i_3_12 = shift_i_map_32;
      6'b100001 : _zz_shift_i_3_12 = shift_i_map_33;
      6'b100010 : _zz_shift_i_3_12 = shift_i_map_34;
      6'b100011 : _zz_shift_i_3_12 = shift_i_map_35;
      6'b100100 : _zz_shift_i_3_12 = shift_i_map_36;
      6'b100101 : _zz_shift_i_3_12 = shift_i_map_37;
      6'b100110 : _zz_shift_i_3_12 = shift_i_map_38;
      6'b100111 : _zz_shift_i_3_12 = shift_i_map_39;
      6'b101000 : _zz_shift_i_3_12 = shift_i_map_40;
      6'b101001 : _zz_shift_i_3_12 = shift_i_map_41;
      6'b101010 : _zz_shift_i_3_12 = shift_i_map_42;
      6'b101011 : _zz_shift_i_3_12 = shift_i_map_43;
      6'b101100 : _zz_shift_i_3_12 = shift_i_map_44;
      6'b101101 : _zz_shift_i_3_12 = shift_i_map_45;
      6'b101110 : _zz_shift_i_3_12 = shift_i_map_46;
      6'b101111 : _zz_shift_i_3_12 = shift_i_map_47;
      6'b110000 : _zz_shift_i_3_12 = shift_i_map_48;
      6'b110001 : _zz_shift_i_3_12 = shift_i_map_49;
      6'b110010 : _zz_shift_i_3_12 = shift_i_map_50;
      6'b110011 : _zz_shift_i_3_12 = shift_i_map_51;
      6'b110100 : _zz_shift_i_3_12 = shift_i_map_52;
      6'b110101 : _zz_shift_i_3_12 = shift_i_map_53;
      6'b110110 : _zz_shift_i_3_12 = shift_i_map_54;
      6'b110111 : _zz_shift_i_3_12 = shift_i_map_55;
      6'b111000 : _zz_shift_i_3_12 = shift_i_map_56;
      6'b111001 : _zz_shift_i_3_12 = shift_i_map_57;
      6'b111010 : _zz_shift_i_3_12 = shift_i_map_58;
      6'b111011 : _zz_shift_i_3_12 = shift_i_map_59;
      6'b111100 : _zz_shift_i_3_12 = shift_i_map_60;
      6'b111101 : _zz_shift_i_3_12 = shift_i_map_61;
      6'b111110 : _zz_shift_i_3_12 = shift_i_map_62;
      default : _zz_shift_i_3_12 = shift_i_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_3_13)
      6'b000000 : _zz_shift_q_3_12 = shift_q_map_0;
      6'b000001 : _zz_shift_q_3_12 = shift_q_map_1;
      6'b000010 : _zz_shift_q_3_12 = shift_q_map_2;
      6'b000011 : _zz_shift_q_3_12 = shift_q_map_3;
      6'b000100 : _zz_shift_q_3_12 = shift_q_map_4;
      6'b000101 : _zz_shift_q_3_12 = shift_q_map_5;
      6'b000110 : _zz_shift_q_3_12 = shift_q_map_6;
      6'b000111 : _zz_shift_q_3_12 = shift_q_map_7;
      6'b001000 : _zz_shift_q_3_12 = shift_q_map_8;
      6'b001001 : _zz_shift_q_3_12 = shift_q_map_9;
      6'b001010 : _zz_shift_q_3_12 = shift_q_map_10;
      6'b001011 : _zz_shift_q_3_12 = shift_q_map_11;
      6'b001100 : _zz_shift_q_3_12 = shift_q_map_12;
      6'b001101 : _zz_shift_q_3_12 = shift_q_map_13;
      6'b001110 : _zz_shift_q_3_12 = shift_q_map_14;
      6'b001111 : _zz_shift_q_3_12 = shift_q_map_15;
      6'b010000 : _zz_shift_q_3_12 = shift_q_map_16;
      6'b010001 : _zz_shift_q_3_12 = shift_q_map_17;
      6'b010010 : _zz_shift_q_3_12 = shift_q_map_18;
      6'b010011 : _zz_shift_q_3_12 = shift_q_map_19;
      6'b010100 : _zz_shift_q_3_12 = shift_q_map_20;
      6'b010101 : _zz_shift_q_3_12 = shift_q_map_21;
      6'b010110 : _zz_shift_q_3_12 = shift_q_map_22;
      6'b010111 : _zz_shift_q_3_12 = shift_q_map_23;
      6'b011000 : _zz_shift_q_3_12 = shift_q_map_24;
      6'b011001 : _zz_shift_q_3_12 = shift_q_map_25;
      6'b011010 : _zz_shift_q_3_12 = shift_q_map_26;
      6'b011011 : _zz_shift_q_3_12 = shift_q_map_27;
      6'b011100 : _zz_shift_q_3_12 = shift_q_map_28;
      6'b011101 : _zz_shift_q_3_12 = shift_q_map_29;
      6'b011110 : _zz_shift_q_3_12 = shift_q_map_30;
      6'b011111 : _zz_shift_q_3_12 = shift_q_map_31;
      6'b100000 : _zz_shift_q_3_12 = shift_q_map_32;
      6'b100001 : _zz_shift_q_3_12 = shift_q_map_33;
      6'b100010 : _zz_shift_q_3_12 = shift_q_map_34;
      6'b100011 : _zz_shift_q_3_12 = shift_q_map_35;
      6'b100100 : _zz_shift_q_3_12 = shift_q_map_36;
      6'b100101 : _zz_shift_q_3_12 = shift_q_map_37;
      6'b100110 : _zz_shift_q_3_12 = shift_q_map_38;
      6'b100111 : _zz_shift_q_3_12 = shift_q_map_39;
      6'b101000 : _zz_shift_q_3_12 = shift_q_map_40;
      6'b101001 : _zz_shift_q_3_12 = shift_q_map_41;
      6'b101010 : _zz_shift_q_3_12 = shift_q_map_42;
      6'b101011 : _zz_shift_q_3_12 = shift_q_map_43;
      6'b101100 : _zz_shift_q_3_12 = shift_q_map_44;
      6'b101101 : _zz_shift_q_3_12 = shift_q_map_45;
      6'b101110 : _zz_shift_q_3_12 = shift_q_map_46;
      6'b101111 : _zz_shift_q_3_12 = shift_q_map_47;
      6'b110000 : _zz_shift_q_3_12 = shift_q_map_48;
      6'b110001 : _zz_shift_q_3_12 = shift_q_map_49;
      6'b110010 : _zz_shift_q_3_12 = shift_q_map_50;
      6'b110011 : _zz_shift_q_3_12 = shift_q_map_51;
      6'b110100 : _zz_shift_q_3_12 = shift_q_map_52;
      6'b110101 : _zz_shift_q_3_12 = shift_q_map_53;
      6'b110110 : _zz_shift_q_3_12 = shift_q_map_54;
      6'b110111 : _zz_shift_q_3_12 = shift_q_map_55;
      6'b111000 : _zz_shift_q_3_12 = shift_q_map_56;
      6'b111001 : _zz_shift_q_3_12 = shift_q_map_57;
      6'b111010 : _zz_shift_q_3_12 = shift_q_map_58;
      6'b111011 : _zz_shift_q_3_12 = shift_q_map_59;
      6'b111100 : _zz_shift_q_3_12 = shift_q_map_60;
      6'b111101 : _zz_shift_q_3_12 = shift_q_map_61;
      6'b111110 : _zz_shift_q_3_12 = shift_q_map_62;
      default : _zz_shift_q_3_12 = shift_q_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_4_13)
      6'b000000 : _zz_shift_i_4_12 = shift_i_map_0;
      6'b000001 : _zz_shift_i_4_12 = shift_i_map_1;
      6'b000010 : _zz_shift_i_4_12 = shift_i_map_2;
      6'b000011 : _zz_shift_i_4_12 = shift_i_map_3;
      6'b000100 : _zz_shift_i_4_12 = shift_i_map_4;
      6'b000101 : _zz_shift_i_4_12 = shift_i_map_5;
      6'b000110 : _zz_shift_i_4_12 = shift_i_map_6;
      6'b000111 : _zz_shift_i_4_12 = shift_i_map_7;
      6'b001000 : _zz_shift_i_4_12 = shift_i_map_8;
      6'b001001 : _zz_shift_i_4_12 = shift_i_map_9;
      6'b001010 : _zz_shift_i_4_12 = shift_i_map_10;
      6'b001011 : _zz_shift_i_4_12 = shift_i_map_11;
      6'b001100 : _zz_shift_i_4_12 = shift_i_map_12;
      6'b001101 : _zz_shift_i_4_12 = shift_i_map_13;
      6'b001110 : _zz_shift_i_4_12 = shift_i_map_14;
      6'b001111 : _zz_shift_i_4_12 = shift_i_map_15;
      6'b010000 : _zz_shift_i_4_12 = shift_i_map_16;
      6'b010001 : _zz_shift_i_4_12 = shift_i_map_17;
      6'b010010 : _zz_shift_i_4_12 = shift_i_map_18;
      6'b010011 : _zz_shift_i_4_12 = shift_i_map_19;
      6'b010100 : _zz_shift_i_4_12 = shift_i_map_20;
      6'b010101 : _zz_shift_i_4_12 = shift_i_map_21;
      6'b010110 : _zz_shift_i_4_12 = shift_i_map_22;
      6'b010111 : _zz_shift_i_4_12 = shift_i_map_23;
      6'b011000 : _zz_shift_i_4_12 = shift_i_map_24;
      6'b011001 : _zz_shift_i_4_12 = shift_i_map_25;
      6'b011010 : _zz_shift_i_4_12 = shift_i_map_26;
      6'b011011 : _zz_shift_i_4_12 = shift_i_map_27;
      6'b011100 : _zz_shift_i_4_12 = shift_i_map_28;
      6'b011101 : _zz_shift_i_4_12 = shift_i_map_29;
      6'b011110 : _zz_shift_i_4_12 = shift_i_map_30;
      6'b011111 : _zz_shift_i_4_12 = shift_i_map_31;
      6'b100000 : _zz_shift_i_4_12 = shift_i_map_32;
      6'b100001 : _zz_shift_i_4_12 = shift_i_map_33;
      6'b100010 : _zz_shift_i_4_12 = shift_i_map_34;
      6'b100011 : _zz_shift_i_4_12 = shift_i_map_35;
      6'b100100 : _zz_shift_i_4_12 = shift_i_map_36;
      6'b100101 : _zz_shift_i_4_12 = shift_i_map_37;
      6'b100110 : _zz_shift_i_4_12 = shift_i_map_38;
      6'b100111 : _zz_shift_i_4_12 = shift_i_map_39;
      6'b101000 : _zz_shift_i_4_12 = shift_i_map_40;
      6'b101001 : _zz_shift_i_4_12 = shift_i_map_41;
      6'b101010 : _zz_shift_i_4_12 = shift_i_map_42;
      6'b101011 : _zz_shift_i_4_12 = shift_i_map_43;
      6'b101100 : _zz_shift_i_4_12 = shift_i_map_44;
      6'b101101 : _zz_shift_i_4_12 = shift_i_map_45;
      6'b101110 : _zz_shift_i_4_12 = shift_i_map_46;
      6'b101111 : _zz_shift_i_4_12 = shift_i_map_47;
      6'b110000 : _zz_shift_i_4_12 = shift_i_map_48;
      6'b110001 : _zz_shift_i_4_12 = shift_i_map_49;
      6'b110010 : _zz_shift_i_4_12 = shift_i_map_50;
      6'b110011 : _zz_shift_i_4_12 = shift_i_map_51;
      6'b110100 : _zz_shift_i_4_12 = shift_i_map_52;
      6'b110101 : _zz_shift_i_4_12 = shift_i_map_53;
      6'b110110 : _zz_shift_i_4_12 = shift_i_map_54;
      6'b110111 : _zz_shift_i_4_12 = shift_i_map_55;
      6'b111000 : _zz_shift_i_4_12 = shift_i_map_56;
      6'b111001 : _zz_shift_i_4_12 = shift_i_map_57;
      6'b111010 : _zz_shift_i_4_12 = shift_i_map_58;
      6'b111011 : _zz_shift_i_4_12 = shift_i_map_59;
      6'b111100 : _zz_shift_i_4_12 = shift_i_map_60;
      6'b111101 : _zz_shift_i_4_12 = shift_i_map_61;
      6'b111110 : _zz_shift_i_4_12 = shift_i_map_62;
      default : _zz_shift_i_4_12 = shift_i_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_4_13)
      6'b000000 : _zz_shift_q_4_12 = shift_q_map_0;
      6'b000001 : _zz_shift_q_4_12 = shift_q_map_1;
      6'b000010 : _zz_shift_q_4_12 = shift_q_map_2;
      6'b000011 : _zz_shift_q_4_12 = shift_q_map_3;
      6'b000100 : _zz_shift_q_4_12 = shift_q_map_4;
      6'b000101 : _zz_shift_q_4_12 = shift_q_map_5;
      6'b000110 : _zz_shift_q_4_12 = shift_q_map_6;
      6'b000111 : _zz_shift_q_4_12 = shift_q_map_7;
      6'b001000 : _zz_shift_q_4_12 = shift_q_map_8;
      6'b001001 : _zz_shift_q_4_12 = shift_q_map_9;
      6'b001010 : _zz_shift_q_4_12 = shift_q_map_10;
      6'b001011 : _zz_shift_q_4_12 = shift_q_map_11;
      6'b001100 : _zz_shift_q_4_12 = shift_q_map_12;
      6'b001101 : _zz_shift_q_4_12 = shift_q_map_13;
      6'b001110 : _zz_shift_q_4_12 = shift_q_map_14;
      6'b001111 : _zz_shift_q_4_12 = shift_q_map_15;
      6'b010000 : _zz_shift_q_4_12 = shift_q_map_16;
      6'b010001 : _zz_shift_q_4_12 = shift_q_map_17;
      6'b010010 : _zz_shift_q_4_12 = shift_q_map_18;
      6'b010011 : _zz_shift_q_4_12 = shift_q_map_19;
      6'b010100 : _zz_shift_q_4_12 = shift_q_map_20;
      6'b010101 : _zz_shift_q_4_12 = shift_q_map_21;
      6'b010110 : _zz_shift_q_4_12 = shift_q_map_22;
      6'b010111 : _zz_shift_q_4_12 = shift_q_map_23;
      6'b011000 : _zz_shift_q_4_12 = shift_q_map_24;
      6'b011001 : _zz_shift_q_4_12 = shift_q_map_25;
      6'b011010 : _zz_shift_q_4_12 = shift_q_map_26;
      6'b011011 : _zz_shift_q_4_12 = shift_q_map_27;
      6'b011100 : _zz_shift_q_4_12 = shift_q_map_28;
      6'b011101 : _zz_shift_q_4_12 = shift_q_map_29;
      6'b011110 : _zz_shift_q_4_12 = shift_q_map_30;
      6'b011111 : _zz_shift_q_4_12 = shift_q_map_31;
      6'b100000 : _zz_shift_q_4_12 = shift_q_map_32;
      6'b100001 : _zz_shift_q_4_12 = shift_q_map_33;
      6'b100010 : _zz_shift_q_4_12 = shift_q_map_34;
      6'b100011 : _zz_shift_q_4_12 = shift_q_map_35;
      6'b100100 : _zz_shift_q_4_12 = shift_q_map_36;
      6'b100101 : _zz_shift_q_4_12 = shift_q_map_37;
      6'b100110 : _zz_shift_q_4_12 = shift_q_map_38;
      6'b100111 : _zz_shift_q_4_12 = shift_q_map_39;
      6'b101000 : _zz_shift_q_4_12 = shift_q_map_40;
      6'b101001 : _zz_shift_q_4_12 = shift_q_map_41;
      6'b101010 : _zz_shift_q_4_12 = shift_q_map_42;
      6'b101011 : _zz_shift_q_4_12 = shift_q_map_43;
      6'b101100 : _zz_shift_q_4_12 = shift_q_map_44;
      6'b101101 : _zz_shift_q_4_12 = shift_q_map_45;
      6'b101110 : _zz_shift_q_4_12 = shift_q_map_46;
      6'b101111 : _zz_shift_q_4_12 = shift_q_map_47;
      6'b110000 : _zz_shift_q_4_12 = shift_q_map_48;
      6'b110001 : _zz_shift_q_4_12 = shift_q_map_49;
      6'b110010 : _zz_shift_q_4_12 = shift_q_map_50;
      6'b110011 : _zz_shift_q_4_12 = shift_q_map_51;
      6'b110100 : _zz_shift_q_4_12 = shift_q_map_52;
      6'b110101 : _zz_shift_q_4_12 = shift_q_map_53;
      6'b110110 : _zz_shift_q_4_12 = shift_q_map_54;
      6'b110111 : _zz_shift_q_4_12 = shift_q_map_55;
      6'b111000 : _zz_shift_q_4_12 = shift_q_map_56;
      6'b111001 : _zz_shift_q_4_12 = shift_q_map_57;
      6'b111010 : _zz_shift_q_4_12 = shift_q_map_58;
      6'b111011 : _zz_shift_q_4_12 = shift_q_map_59;
      6'b111100 : _zz_shift_q_4_12 = shift_q_map_60;
      6'b111101 : _zz_shift_q_4_12 = shift_q_map_61;
      6'b111110 : _zz_shift_q_4_12 = shift_q_map_62;
      default : _zz_shift_q_4_12 = shift_q_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_5_13)
      6'b000000 : _zz_shift_i_5_12 = shift_i_map_0;
      6'b000001 : _zz_shift_i_5_12 = shift_i_map_1;
      6'b000010 : _zz_shift_i_5_12 = shift_i_map_2;
      6'b000011 : _zz_shift_i_5_12 = shift_i_map_3;
      6'b000100 : _zz_shift_i_5_12 = shift_i_map_4;
      6'b000101 : _zz_shift_i_5_12 = shift_i_map_5;
      6'b000110 : _zz_shift_i_5_12 = shift_i_map_6;
      6'b000111 : _zz_shift_i_5_12 = shift_i_map_7;
      6'b001000 : _zz_shift_i_5_12 = shift_i_map_8;
      6'b001001 : _zz_shift_i_5_12 = shift_i_map_9;
      6'b001010 : _zz_shift_i_5_12 = shift_i_map_10;
      6'b001011 : _zz_shift_i_5_12 = shift_i_map_11;
      6'b001100 : _zz_shift_i_5_12 = shift_i_map_12;
      6'b001101 : _zz_shift_i_5_12 = shift_i_map_13;
      6'b001110 : _zz_shift_i_5_12 = shift_i_map_14;
      6'b001111 : _zz_shift_i_5_12 = shift_i_map_15;
      6'b010000 : _zz_shift_i_5_12 = shift_i_map_16;
      6'b010001 : _zz_shift_i_5_12 = shift_i_map_17;
      6'b010010 : _zz_shift_i_5_12 = shift_i_map_18;
      6'b010011 : _zz_shift_i_5_12 = shift_i_map_19;
      6'b010100 : _zz_shift_i_5_12 = shift_i_map_20;
      6'b010101 : _zz_shift_i_5_12 = shift_i_map_21;
      6'b010110 : _zz_shift_i_5_12 = shift_i_map_22;
      6'b010111 : _zz_shift_i_5_12 = shift_i_map_23;
      6'b011000 : _zz_shift_i_5_12 = shift_i_map_24;
      6'b011001 : _zz_shift_i_5_12 = shift_i_map_25;
      6'b011010 : _zz_shift_i_5_12 = shift_i_map_26;
      6'b011011 : _zz_shift_i_5_12 = shift_i_map_27;
      6'b011100 : _zz_shift_i_5_12 = shift_i_map_28;
      6'b011101 : _zz_shift_i_5_12 = shift_i_map_29;
      6'b011110 : _zz_shift_i_5_12 = shift_i_map_30;
      6'b011111 : _zz_shift_i_5_12 = shift_i_map_31;
      6'b100000 : _zz_shift_i_5_12 = shift_i_map_32;
      6'b100001 : _zz_shift_i_5_12 = shift_i_map_33;
      6'b100010 : _zz_shift_i_5_12 = shift_i_map_34;
      6'b100011 : _zz_shift_i_5_12 = shift_i_map_35;
      6'b100100 : _zz_shift_i_5_12 = shift_i_map_36;
      6'b100101 : _zz_shift_i_5_12 = shift_i_map_37;
      6'b100110 : _zz_shift_i_5_12 = shift_i_map_38;
      6'b100111 : _zz_shift_i_5_12 = shift_i_map_39;
      6'b101000 : _zz_shift_i_5_12 = shift_i_map_40;
      6'b101001 : _zz_shift_i_5_12 = shift_i_map_41;
      6'b101010 : _zz_shift_i_5_12 = shift_i_map_42;
      6'b101011 : _zz_shift_i_5_12 = shift_i_map_43;
      6'b101100 : _zz_shift_i_5_12 = shift_i_map_44;
      6'b101101 : _zz_shift_i_5_12 = shift_i_map_45;
      6'b101110 : _zz_shift_i_5_12 = shift_i_map_46;
      6'b101111 : _zz_shift_i_5_12 = shift_i_map_47;
      6'b110000 : _zz_shift_i_5_12 = shift_i_map_48;
      6'b110001 : _zz_shift_i_5_12 = shift_i_map_49;
      6'b110010 : _zz_shift_i_5_12 = shift_i_map_50;
      6'b110011 : _zz_shift_i_5_12 = shift_i_map_51;
      6'b110100 : _zz_shift_i_5_12 = shift_i_map_52;
      6'b110101 : _zz_shift_i_5_12 = shift_i_map_53;
      6'b110110 : _zz_shift_i_5_12 = shift_i_map_54;
      6'b110111 : _zz_shift_i_5_12 = shift_i_map_55;
      6'b111000 : _zz_shift_i_5_12 = shift_i_map_56;
      6'b111001 : _zz_shift_i_5_12 = shift_i_map_57;
      6'b111010 : _zz_shift_i_5_12 = shift_i_map_58;
      6'b111011 : _zz_shift_i_5_12 = shift_i_map_59;
      6'b111100 : _zz_shift_i_5_12 = shift_i_map_60;
      6'b111101 : _zz_shift_i_5_12 = shift_i_map_61;
      6'b111110 : _zz_shift_i_5_12 = shift_i_map_62;
      default : _zz_shift_i_5_12 = shift_i_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_5_13)
      6'b000000 : _zz_shift_q_5_12 = shift_q_map_0;
      6'b000001 : _zz_shift_q_5_12 = shift_q_map_1;
      6'b000010 : _zz_shift_q_5_12 = shift_q_map_2;
      6'b000011 : _zz_shift_q_5_12 = shift_q_map_3;
      6'b000100 : _zz_shift_q_5_12 = shift_q_map_4;
      6'b000101 : _zz_shift_q_5_12 = shift_q_map_5;
      6'b000110 : _zz_shift_q_5_12 = shift_q_map_6;
      6'b000111 : _zz_shift_q_5_12 = shift_q_map_7;
      6'b001000 : _zz_shift_q_5_12 = shift_q_map_8;
      6'b001001 : _zz_shift_q_5_12 = shift_q_map_9;
      6'b001010 : _zz_shift_q_5_12 = shift_q_map_10;
      6'b001011 : _zz_shift_q_5_12 = shift_q_map_11;
      6'b001100 : _zz_shift_q_5_12 = shift_q_map_12;
      6'b001101 : _zz_shift_q_5_12 = shift_q_map_13;
      6'b001110 : _zz_shift_q_5_12 = shift_q_map_14;
      6'b001111 : _zz_shift_q_5_12 = shift_q_map_15;
      6'b010000 : _zz_shift_q_5_12 = shift_q_map_16;
      6'b010001 : _zz_shift_q_5_12 = shift_q_map_17;
      6'b010010 : _zz_shift_q_5_12 = shift_q_map_18;
      6'b010011 : _zz_shift_q_5_12 = shift_q_map_19;
      6'b010100 : _zz_shift_q_5_12 = shift_q_map_20;
      6'b010101 : _zz_shift_q_5_12 = shift_q_map_21;
      6'b010110 : _zz_shift_q_5_12 = shift_q_map_22;
      6'b010111 : _zz_shift_q_5_12 = shift_q_map_23;
      6'b011000 : _zz_shift_q_5_12 = shift_q_map_24;
      6'b011001 : _zz_shift_q_5_12 = shift_q_map_25;
      6'b011010 : _zz_shift_q_5_12 = shift_q_map_26;
      6'b011011 : _zz_shift_q_5_12 = shift_q_map_27;
      6'b011100 : _zz_shift_q_5_12 = shift_q_map_28;
      6'b011101 : _zz_shift_q_5_12 = shift_q_map_29;
      6'b011110 : _zz_shift_q_5_12 = shift_q_map_30;
      6'b011111 : _zz_shift_q_5_12 = shift_q_map_31;
      6'b100000 : _zz_shift_q_5_12 = shift_q_map_32;
      6'b100001 : _zz_shift_q_5_12 = shift_q_map_33;
      6'b100010 : _zz_shift_q_5_12 = shift_q_map_34;
      6'b100011 : _zz_shift_q_5_12 = shift_q_map_35;
      6'b100100 : _zz_shift_q_5_12 = shift_q_map_36;
      6'b100101 : _zz_shift_q_5_12 = shift_q_map_37;
      6'b100110 : _zz_shift_q_5_12 = shift_q_map_38;
      6'b100111 : _zz_shift_q_5_12 = shift_q_map_39;
      6'b101000 : _zz_shift_q_5_12 = shift_q_map_40;
      6'b101001 : _zz_shift_q_5_12 = shift_q_map_41;
      6'b101010 : _zz_shift_q_5_12 = shift_q_map_42;
      6'b101011 : _zz_shift_q_5_12 = shift_q_map_43;
      6'b101100 : _zz_shift_q_5_12 = shift_q_map_44;
      6'b101101 : _zz_shift_q_5_12 = shift_q_map_45;
      6'b101110 : _zz_shift_q_5_12 = shift_q_map_46;
      6'b101111 : _zz_shift_q_5_12 = shift_q_map_47;
      6'b110000 : _zz_shift_q_5_12 = shift_q_map_48;
      6'b110001 : _zz_shift_q_5_12 = shift_q_map_49;
      6'b110010 : _zz_shift_q_5_12 = shift_q_map_50;
      6'b110011 : _zz_shift_q_5_12 = shift_q_map_51;
      6'b110100 : _zz_shift_q_5_12 = shift_q_map_52;
      6'b110101 : _zz_shift_q_5_12 = shift_q_map_53;
      6'b110110 : _zz_shift_q_5_12 = shift_q_map_54;
      6'b110111 : _zz_shift_q_5_12 = shift_q_map_55;
      6'b111000 : _zz_shift_q_5_12 = shift_q_map_56;
      6'b111001 : _zz_shift_q_5_12 = shift_q_map_57;
      6'b111010 : _zz_shift_q_5_12 = shift_q_map_58;
      6'b111011 : _zz_shift_q_5_12 = shift_q_map_59;
      6'b111100 : _zz_shift_q_5_12 = shift_q_map_60;
      6'b111101 : _zz_shift_q_5_12 = shift_q_map_61;
      6'b111110 : _zz_shift_q_5_12 = shift_q_map_62;
      default : _zz_shift_q_5_12 = shift_q_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_6_13)
      6'b000000 : _zz_shift_i_6_12 = shift_i_map_0;
      6'b000001 : _zz_shift_i_6_12 = shift_i_map_1;
      6'b000010 : _zz_shift_i_6_12 = shift_i_map_2;
      6'b000011 : _zz_shift_i_6_12 = shift_i_map_3;
      6'b000100 : _zz_shift_i_6_12 = shift_i_map_4;
      6'b000101 : _zz_shift_i_6_12 = shift_i_map_5;
      6'b000110 : _zz_shift_i_6_12 = shift_i_map_6;
      6'b000111 : _zz_shift_i_6_12 = shift_i_map_7;
      6'b001000 : _zz_shift_i_6_12 = shift_i_map_8;
      6'b001001 : _zz_shift_i_6_12 = shift_i_map_9;
      6'b001010 : _zz_shift_i_6_12 = shift_i_map_10;
      6'b001011 : _zz_shift_i_6_12 = shift_i_map_11;
      6'b001100 : _zz_shift_i_6_12 = shift_i_map_12;
      6'b001101 : _zz_shift_i_6_12 = shift_i_map_13;
      6'b001110 : _zz_shift_i_6_12 = shift_i_map_14;
      6'b001111 : _zz_shift_i_6_12 = shift_i_map_15;
      6'b010000 : _zz_shift_i_6_12 = shift_i_map_16;
      6'b010001 : _zz_shift_i_6_12 = shift_i_map_17;
      6'b010010 : _zz_shift_i_6_12 = shift_i_map_18;
      6'b010011 : _zz_shift_i_6_12 = shift_i_map_19;
      6'b010100 : _zz_shift_i_6_12 = shift_i_map_20;
      6'b010101 : _zz_shift_i_6_12 = shift_i_map_21;
      6'b010110 : _zz_shift_i_6_12 = shift_i_map_22;
      6'b010111 : _zz_shift_i_6_12 = shift_i_map_23;
      6'b011000 : _zz_shift_i_6_12 = shift_i_map_24;
      6'b011001 : _zz_shift_i_6_12 = shift_i_map_25;
      6'b011010 : _zz_shift_i_6_12 = shift_i_map_26;
      6'b011011 : _zz_shift_i_6_12 = shift_i_map_27;
      6'b011100 : _zz_shift_i_6_12 = shift_i_map_28;
      6'b011101 : _zz_shift_i_6_12 = shift_i_map_29;
      6'b011110 : _zz_shift_i_6_12 = shift_i_map_30;
      6'b011111 : _zz_shift_i_6_12 = shift_i_map_31;
      6'b100000 : _zz_shift_i_6_12 = shift_i_map_32;
      6'b100001 : _zz_shift_i_6_12 = shift_i_map_33;
      6'b100010 : _zz_shift_i_6_12 = shift_i_map_34;
      6'b100011 : _zz_shift_i_6_12 = shift_i_map_35;
      6'b100100 : _zz_shift_i_6_12 = shift_i_map_36;
      6'b100101 : _zz_shift_i_6_12 = shift_i_map_37;
      6'b100110 : _zz_shift_i_6_12 = shift_i_map_38;
      6'b100111 : _zz_shift_i_6_12 = shift_i_map_39;
      6'b101000 : _zz_shift_i_6_12 = shift_i_map_40;
      6'b101001 : _zz_shift_i_6_12 = shift_i_map_41;
      6'b101010 : _zz_shift_i_6_12 = shift_i_map_42;
      6'b101011 : _zz_shift_i_6_12 = shift_i_map_43;
      6'b101100 : _zz_shift_i_6_12 = shift_i_map_44;
      6'b101101 : _zz_shift_i_6_12 = shift_i_map_45;
      6'b101110 : _zz_shift_i_6_12 = shift_i_map_46;
      6'b101111 : _zz_shift_i_6_12 = shift_i_map_47;
      6'b110000 : _zz_shift_i_6_12 = shift_i_map_48;
      6'b110001 : _zz_shift_i_6_12 = shift_i_map_49;
      6'b110010 : _zz_shift_i_6_12 = shift_i_map_50;
      6'b110011 : _zz_shift_i_6_12 = shift_i_map_51;
      6'b110100 : _zz_shift_i_6_12 = shift_i_map_52;
      6'b110101 : _zz_shift_i_6_12 = shift_i_map_53;
      6'b110110 : _zz_shift_i_6_12 = shift_i_map_54;
      6'b110111 : _zz_shift_i_6_12 = shift_i_map_55;
      6'b111000 : _zz_shift_i_6_12 = shift_i_map_56;
      6'b111001 : _zz_shift_i_6_12 = shift_i_map_57;
      6'b111010 : _zz_shift_i_6_12 = shift_i_map_58;
      6'b111011 : _zz_shift_i_6_12 = shift_i_map_59;
      6'b111100 : _zz_shift_i_6_12 = shift_i_map_60;
      6'b111101 : _zz_shift_i_6_12 = shift_i_map_61;
      6'b111110 : _zz_shift_i_6_12 = shift_i_map_62;
      default : _zz_shift_i_6_12 = shift_i_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_6_13)
      6'b000000 : _zz_shift_q_6_12 = shift_q_map_0;
      6'b000001 : _zz_shift_q_6_12 = shift_q_map_1;
      6'b000010 : _zz_shift_q_6_12 = shift_q_map_2;
      6'b000011 : _zz_shift_q_6_12 = shift_q_map_3;
      6'b000100 : _zz_shift_q_6_12 = shift_q_map_4;
      6'b000101 : _zz_shift_q_6_12 = shift_q_map_5;
      6'b000110 : _zz_shift_q_6_12 = shift_q_map_6;
      6'b000111 : _zz_shift_q_6_12 = shift_q_map_7;
      6'b001000 : _zz_shift_q_6_12 = shift_q_map_8;
      6'b001001 : _zz_shift_q_6_12 = shift_q_map_9;
      6'b001010 : _zz_shift_q_6_12 = shift_q_map_10;
      6'b001011 : _zz_shift_q_6_12 = shift_q_map_11;
      6'b001100 : _zz_shift_q_6_12 = shift_q_map_12;
      6'b001101 : _zz_shift_q_6_12 = shift_q_map_13;
      6'b001110 : _zz_shift_q_6_12 = shift_q_map_14;
      6'b001111 : _zz_shift_q_6_12 = shift_q_map_15;
      6'b010000 : _zz_shift_q_6_12 = shift_q_map_16;
      6'b010001 : _zz_shift_q_6_12 = shift_q_map_17;
      6'b010010 : _zz_shift_q_6_12 = shift_q_map_18;
      6'b010011 : _zz_shift_q_6_12 = shift_q_map_19;
      6'b010100 : _zz_shift_q_6_12 = shift_q_map_20;
      6'b010101 : _zz_shift_q_6_12 = shift_q_map_21;
      6'b010110 : _zz_shift_q_6_12 = shift_q_map_22;
      6'b010111 : _zz_shift_q_6_12 = shift_q_map_23;
      6'b011000 : _zz_shift_q_6_12 = shift_q_map_24;
      6'b011001 : _zz_shift_q_6_12 = shift_q_map_25;
      6'b011010 : _zz_shift_q_6_12 = shift_q_map_26;
      6'b011011 : _zz_shift_q_6_12 = shift_q_map_27;
      6'b011100 : _zz_shift_q_6_12 = shift_q_map_28;
      6'b011101 : _zz_shift_q_6_12 = shift_q_map_29;
      6'b011110 : _zz_shift_q_6_12 = shift_q_map_30;
      6'b011111 : _zz_shift_q_6_12 = shift_q_map_31;
      6'b100000 : _zz_shift_q_6_12 = shift_q_map_32;
      6'b100001 : _zz_shift_q_6_12 = shift_q_map_33;
      6'b100010 : _zz_shift_q_6_12 = shift_q_map_34;
      6'b100011 : _zz_shift_q_6_12 = shift_q_map_35;
      6'b100100 : _zz_shift_q_6_12 = shift_q_map_36;
      6'b100101 : _zz_shift_q_6_12 = shift_q_map_37;
      6'b100110 : _zz_shift_q_6_12 = shift_q_map_38;
      6'b100111 : _zz_shift_q_6_12 = shift_q_map_39;
      6'b101000 : _zz_shift_q_6_12 = shift_q_map_40;
      6'b101001 : _zz_shift_q_6_12 = shift_q_map_41;
      6'b101010 : _zz_shift_q_6_12 = shift_q_map_42;
      6'b101011 : _zz_shift_q_6_12 = shift_q_map_43;
      6'b101100 : _zz_shift_q_6_12 = shift_q_map_44;
      6'b101101 : _zz_shift_q_6_12 = shift_q_map_45;
      6'b101110 : _zz_shift_q_6_12 = shift_q_map_46;
      6'b101111 : _zz_shift_q_6_12 = shift_q_map_47;
      6'b110000 : _zz_shift_q_6_12 = shift_q_map_48;
      6'b110001 : _zz_shift_q_6_12 = shift_q_map_49;
      6'b110010 : _zz_shift_q_6_12 = shift_q_map_50;
      6'b110011 : _zz_shift_q_6_12 = shift_q_map_51;
      6'b110100 : _zz_shift_q_6_12 = shift_q_map_52;
      6'b110101 : _zz_shift_q_6_12 = shift_q_map_53;
      6'b110110 : _zz_shift_q_6_12 = shift_q_map_54;
      6'b110111 : _zz_shift_q_6_12 = shift_q_map_55;
      6'b111000 : _zz_shift_q_6_12 = shift_q_map_56;
      6'b111001 : _zz_shift_q_6_12 = shift_q_map_57;
      6'b111010 : _zz_shift_q_6_12 = shift_q_map_58;
      6'b111011 : _zz_shift_q_6_12 = shift_q_map_59;
      6'b111100 : _zz_shift_q_6_12 = shift_q_map_60;
      6'b111101 : _zz_shift_q_6_12 = shift_q_map_61;
      6'b111110 : _zz_shift_q_6_12 = shift_q_map_62;
      default : _zz_shift_q_6_12 = shift_q_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_7_13)
      6'b000000 : _zz_shift_i_7_12 = shift_i_map_0;
      6'b000001 : _zz_shift_i_7_12 = shift_i_map_1;
      6'b000010 : _zz_shift_i_7_12 = shift_i_map_2;
      6'b000011 : _zz_shift_i_7_12 = shift_i_map_3;
      6'b000100 : _zz_shift_i_7_12 = shift_i_map_4;
      6'b000101 : _zz_shift_i_7_12 = shift_i_map_5;
      6'b000110 : _zz_shift_i_7_12 = shift_i_map_6;
      6'b000111 : _zz_shift_i_7_12 = shift_i_map_7;
      6'b001000 : _zz_shift_i_7_12 = shift_i_map_8;
      6'b001001 : _zz_shift_i_7_12 = shift_i_map_9;
      6'b001010 : _zz_shift_i_7_12 = shift_i_map_10;
      6'b001011 : _zz_shift_i_7_12 = shift_i_map_11;
      6'b001100 : _zz_shift_i_7_12 = shift_i_map_12;
      6'b001101 : _zz_shift_i_7_12 = shift_i_map_13;
      6'b001110 : _zz_shift_i_7_12 = shift_i_map_14;
      6'b001111 : _zz_shift_i_7_12 = shift_i_map_15;
      6'b010000 : _zz_shift_i_7_12 = shift_i_map_16;
      6'b010001 : _zz_shift_i_7_12 = shift_i_map_17;
      6'b010010 : _zz_shift_i_7_12 = shift_i_map_18;
      6'b010011 : _zz_shift_i_7_12 = shift_i_map_19;
      6'b010100 : _zz_shift_i_7_12 = shift_i_map_20;
      6'b010101 : _zz_shift_i_7_12 = shift_i_map_21;
      6'b010110 : _zz_shift_i_7_12 = shift_i_map_22;
      6'b010111 : _zz_shift_i_7_12 = shift_i_map_23;
      6'b011000 : _zz_shift_i_7_12 = shift_i_map_24;
      6'b011001 : _zz_shift_i_7_12 = shift_i_map_25;
      6'b011010 : _zz_shift_i_7_12 = shift_i_map_26;
      6'b011011 : _zz_shift_i_7_12 = shift_i_map_27;
      6'b011100 : _zz_shift_i_7_12 = shift_i_map_28;
      6'b011101 : _zz_shift_i_7_12 = shift_i_map_29;
      6'b011110 : _zz_shift_i_7_12 = shift_i_map_30;
      6'b011111 : _zz_shift_i_7_12 = shift_i_map_31;
      6'b100000 : _zz_shift_i_7_12 = shift_i_map_32;
      6'b100001 : _zz_shift_i_7_12 = shift_i_map_33;
      6'b100010 : _zz_shift_i_7_12 = shift_i_map_34;
      6'b100011 : _zz_shift_i_7_12 = shift_i_map_35;
      6'b100100 : _zz_shift_i_7_12 = shift_i_map_36;
      6'b100101 : _zz_shift_i_7_12 = shift_i_map_37;
      6'b100110 : _zz_shift_i_7_12 = shift_i_map_38;
      6'b100111 : _zz_shift_i_7_12 = shift_i_map_39;
      6'b101000 : _zz_shift_i_7_12 = shift_i_map_40;
      6'b101001 : _zz_shift_i_7_12 = shift_i_map_41;
      6'b101010 : _zz_shift_i_7_12 = shift_i_map_42;
      6'b101011 : _zz_shift_i_7_12 = shift_i_map_43;
      6'b101100 : _zz_shift_i_7_12 = shift_i_map_44;
      6'b101101 : _zz_shift_i_7_12 = shift_i_map_45;
      6'b101110 : _zz_shift_i_7_12 = shift_i_map_46;
      6'b101111 : _zz_shift_i_7_12 = shift_i_map_47;
      6'b110000 : _zz_shift_i_7_12 = shift_i_map_48;
      6'b110001 : _zz_shift_i_7_12 = shift_i_map_49;
      6'b110010 : _zz_shift_i_7_12 = shift_i_map_50;
      6'b110011 : _zz_shift_i_7_12 = shift_i_map_51;
      6'b110100 : _zz_shift_i_7_12 = shift_i_map_52;
      6'b110101 : _zz_shift_i_7_12 = shift_i_map_53;
      6'b110110 : _zz_shift_i_7_12 = shift_i_map_54;
      6'b110111 : _zz_shift_i_7_12 = shift_i_map_55;
      6'b111000 : _zz_shift_i_7_12 = shift_i_map_56;
      6'b111001 : _zz_shift_i_7_12 = shift_i_map_57;
      6'b111010 : _zz_shift_i_7_12 = shift_i_map_58;
      6'b111011 : _zz_shift_i_7_12 = shift_i_map_59;
      6'b111100 : _zz_shift_i_7_12 = shift_i_map_60;
      6'b111101 : _zz_shift_i_7_12 = shift_i_map_61;
      6'b111110 : _zz_shift_i_7_12 = shift_i_map_62;
      default : _zz_shift_i_7_12 = shift_i_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_7_13)
      6'b000000 : _zz_shift_q_7_12 = shift_q_map_0;
      6'b000001 : _zz_shift_q_7_12 = shift_q_map_1;
      6'b000010 : _zz_shift_q_7_12 = shift_q_map_2;
      6'b000011 : _zz_shift_q_7_12 = shift_q_map_3;
      6'b000100 : _zz_shift_q_7_12 = shift_q_map_4;
      6'b000101 : _zz_shift_q_7_12 = shift_q_map_5;
      6'b000110 : _zz_shift_q_7_12 = shift_q_map_6;
      6'b000111 : _zz_shift_q_7_12 = shift_q_map_7;
      6'b001000 : _zz_shift_q_7_12 = shift_q_map_8;
      6'b001001 : _zz_shift_q_7_12 = shift_q_map_9;
      6'b001010 : _zz_shift_q_7_12 = shift_q_map_10;
      6'b001011 : _zz_shift_q_7_12 = shift_q_map_11;
      6'b001100 : _zz_shift_q_7_12 = shift_q_map_12;
      6'b001101 : _zz_shift_q_7_12 = shift_q_map_13;
      6'b001110 : _zz_shift_q_7_12 = shift_q_map_14;
      6'b001111 : _zz_shift_q_7_12 = shift_q_map_15;
      6'b010000 : _zz_shift_q_7_12 = shift_q_map_16;
      6'b010001 : _zz_shift_q_7_12 = shift_q_map_17;
      6'b010010 : _zz_shift_q_7_12 = shift_q_map_18;
      6'b010011 : _zz_shift_q_7_12 = shift_q_map_19;
      6'b010100 : _zz_shift_q_7_12 = shift_q_map_20;
      6'b010101 : _zz_shift_q_7_12 = shift_q_map_21;
      6'b010110 : _zz_shift_q_7_12 = shift_q_map_22;
      6'b010111 : _zz_shift_q_7_12 = shift_q_map_23;
      6'b011000 : _zz_shift_q_7_12 = shift_q_map_24;
      6'b011001 : _zz_shift_q_7_12 = shift_q_map_25;
      6'b011010 : _zz_shift_q_7_12 = shift_q_map_26;
      6'b011011 : _zz_shift_q_7_12 = shift_q_map_27;
      6'b011100 : _zz_shift_q_7_12 = shift_q_map_28;
      6'b011101 : _zz_shift_q_7_12 = shift_q_map_29;
      6'b011110 : _zz_shift_q_7_12 = shift_q_map_30;
      6'b011111 : _zz_shift_q_7_12 = shift_q_map_31;
      6'b100000 : _zz_shift_q_7_12 = shift_q_map_32;
      6'b100001 : _zz_shift_q_7_12 = shift_q_map_33;
      6'b100010 : _zz_shift_q_7_12 = shift_q_map_34;
      6'b100011 : _zz_shift_q_7_12 = shift_q_map_35;
      6'b100100 : _zz_shift_q_7_12 = shift_q_map_36;
      6'b100101 : _zz_shift_q_7_12 = shift_q_map_37;
      6'b100110 : _zz_shift_q_7_12 = shift_q_map_38;
      6'b100111 : _zz_shift_q_7_12 = shift_q_map_39;
      6'b101000 : _zz_shift_q_7_12 = shift_q_map_40;
      6'b101001 : _zz_shift_q_7_12 = shift_q_map_41;
      6'b101010 : _zz_shift_q_7_12 = shift_q_map_42;
      6'b101011 : _zz_shift_q_7_12 = shift_q_map_43;
      6'b101100 : _zz_shift_q_7_12 = shift_q_map_44;
      6'b101101 : _zz_shift_q_7_12 = shift_q_map_45;
      6'b101110 : _zz_shift_q_7_12 = shift_q_map_46;
      6'b101111 : _zz_shift_q_7_12 = shift_q_map_47;
      6'b110000 : _zz_shift_q_7_12 = shift_q_map_48;
      6'b110001 : _zz_shift_q_7_12 = shift_q_map_49;
      6'b110010 : _zz_shift_q_7_12 = shift_q_map_50;
      6'b110011 : _zz_shift_q_7_12 = shift_q_map_51;
      6'b110100 : _zz_shift_q_7_12 = shift_q_map_52;
      6'b110101 : _zz_shift_q_7_12 = shift_q_map_53;
      6'b110110 : _zz_shift_q_7_12 = shift_q_map_54;
      6'b110111 : _zz_shift_q_7_12 = shift_q_map_55;
      6'b111000 : _zz_shift_q_7_12 = shift_q_map_56;
      6'b111001 : _zz_shift_q_7_12 = shift_q_map_57;
      6'b111010 : _zz_shift_q_7_12 = shift_q_map_58;
      6'b111011 : _zz_shift_q_7_12 = shift_q_map_59;
      6'b111100 : _zz_shift_q_7_12 = shift_q_map_60;
      6'b111101 : _zz_shift_q_7_12 = shift_q_map_61;
      6'b111110 : _zz_shift_q_7_12 = shift_q_map_62;
      default : _zz_shift_q_7_12 = shift_q_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_0_15)
      6'b000000 : _zz_shift_i_0_14 = shift_i_map_0;
      6'b000001 : _zz_shift_i_0_14 = shift_i_map_1;
      6'b000010 : _zz_shift_i_0_14 = shift_i_map_2;
      6'b000011 : _zz_shift_i_0_14 = shift_i_map_3;
      6'b000100 : _zz_shift_i_0_14 = shift_i_map_4;
      6'b000101 : _zz_shift_i_0_14 = shift_i_map_5;
      6'b000110 : _zz_shift_i_0_14 = shift_i_map_6;
      6'b000111 : _zz_shift_i_0_14 = shift_i_map_7;
      6'b001000 : _zz_shift_i_0_14 = shift_i_map_8;
      6'b001001 : _zz_shift_i_0_14 = shift_i_map_9;
      6'b001010 : _zz_shift_i_0_14 = shift_i_map_10;
      6'b001011 : _zz_shift_i_0_14 = shift_i_map_11;
      6'b001100 : _zz_shift_i_0_14 = shift_i_map_12;
      6'b001101 : _zz_shift_i_0_14 = shift_i_map_13;
      6'b001110 : _zz_shift_i_0_14 = shift_i_map_14;
      6'b001111 : _zz_shift_i_0_14 = shift_i_map_15;
      6'b010000 : _zz_shift_i_0_14 = shift_i_map_16;
      6'b010001 : _zz_shift_i_0_14 = shift_i_map_17;
      6'b010010 : _zz_shift_i_0_14 = shift_i_map_18;
      6'b010011 : _zz_shift_i_0_14 = shift_i_map_19;
      6'b010100 : _zz_shift_i_0_14 = shift_i_map_20;
      6'b010101 : _zz_shift_i_0_14 = shift_i_map_21;
      6'b010110 : _zz_shift_i_0_14 = shift_i_map_22;
      6'b010111 : _zz_shift_i_0_14 = shift_i_map_23;
      6'b011000 : _zz_shift_i_0_14 = shift_i_map_24;
      6'b011001 : _zz_shift_i_0_14 = shift_i_map_25;
      6'b011010 : _zz_shift_i_0_14 = shift_i_map_26;
      6'b011011 : _zz_shift_i_0_14 = shift_i_map_27;
      6'b011100 : _zz_shift_i_0_14 = shift_i_map_28;
      6'b011101 : _zz_shift_i_0_14 = shift_i_map_29;
      6'b011110 : _zz_shift_i_0_14 = shift_i_map_30;
      6'b011111 : _zz_shift_i_0_14 = shift_i_map_31;
      6'b100000 : _zz_shift_i_0_14 = shift_i_map_32;
      6'b100001 : _zz_shift_i_0_14 = shift_i_map_33;
      6'b100010 : _zz_shift_i_0_14 = shift_i_map_34;
      6'b100011 : _zz_shift_i_0_14 = shift_i_map_35;
      6'b100100 : _zz_shift_i_0_14 = shift_i_map_36;
      6'b100101 : _zz_shift_i_0_14 = shift_i_map_37;
      6'b100110 : _zz_shift_i_0_14 = shift_i_map_38;
      6'b100111 : _zz_shift_i_0_14 = shift_i_map_39;
      6'b101000 : _zz_shift_i_0_14 = shift_i_map_40;
      6'b101001 : _zz_shift_i_0_14 = shift_i_map_41;
      6'b101010 : _zz_shift_i_0_14 = shift_i_map_42;
      6'b101011 : _zz_shift_i_0_14 = shift_i_map_43;
      6'b101100 : _zz_shift_i_0_14 = shift_i_map_44;
      6'b101101 : _zz_shift_i_0_14 = shift_i_map_45;
      6'b101110 : _zz_shift_i_0_14 = shift_i_map_46;
      6'b101111 : _zz_shift_i_0_14 = shift_i_map_47;
      6'b110000 : _zz_shift_i_0_14 = shift_i_map_48;
      6'b110001 : _zz_shift_i_0_14 = shift_i_map_49;
      6'b110010 : _zz_shift_i_0_14 = shift_i_map_50;
      6'b110011 : _zz_shift_i_0_14 = shift_i_map_51;
      6'b110100 : _zz_shift_i_0_14 = shift_i_map_52;
      6'b110101 : _zz_shift_i_0_14 = shift_i_map_53;
      6'b110110 : _zz_shift_i_0_14 = shift_i_map_54;
      6'b110111 : _zz_shift_i_0_14 = shift_i_map_55;
      6'b111000 : _zz_shift_i_0_14 = shift_i_map_56;
      6'b111001 : _zz_shift_i_0_14 = shift_i_map_57;
      6'b111010 : _zz_shift_i_0_14 = shift_i_map_58;
      6'b111011 : _zz_shift_i_0_14 = shift_i_map_59;
      6'b111100 : _zz_shift_i_0_14 = shift_i_map_60;
      6'b111101 : _zz_shift_i_0_14 = shift_i_map_61;
      6'b111110 : _zz_shift_i_0_14 = shift_i_map_62;
      default : _zz_shift_i_0_14 = shift_i_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_0_15)
      6'b000000 : _zz_shift_q_0_14 = shift_q_map_0;
      6'b000001 : _zz_shift_q_0_14 = shift_q_map_1;
      6'b000010 : _zz_shift_q_0_14 = shift_q_map_2;
      6'b000011 : _zz_shift_q_0_14 = shift_q_map_3;
      6'b000100 : _zz_shift_q_0_14 = shift_q_map_4;
      6'b000101 : _zz_shift_q_0_14 = shift_q_map_5;
      6'b000110 : _zz_shift_q_0_14 = shift_q_map_6;
      6'b000111 : _zz_shift_q_0_14 = shift_q_map_7;
      6'b001000 : _zz_shift_q_0_14 = shift_q_map_8;
      6'b001001 : _zz_shift_q_0_14 = shift_q_map_9;
      6'b001010 : _zz_shift_q_0_14 = shift_q_map_10;
      6'b001011 : _zz_shift_q_0_14 = shift_q_map_11;
      6'b001100 : _zz_shift_q_0_14 = shift_q_map_12;
      6'b001101 : _zz_shift_q_0_14 = shift_q_map_13;
      6'b001110 : _zz_shift_q_0_14 = shift_q_map_14;
      6'b001111 : _zz_shift_q_0_14 = shift_q_map_15;
      6'b010000 : _zz_shift_q_0_14 = shift_q_map_16;
      6'b010001 : _zz_shift_q_0_14 = shift_q_map_17;
      6'b010010 : _zz_shift_q_0_14 = shift_q_map_18;
      6'b010011 : _zz_shift_q_0_14 = shift_q_map_19;
      6'b010100 : _zz_shift_q_0_14 = shift_q_map_20;
      6'b010101 : _zz_shift_q_0_14 = shift_q_map_21;
      6'b010110 : _zz_shift_q_0_14 = shift_q_map_22;
      6'b010111 : _zz_shift_q_0_14 = shift_q_map_23;
      6'b011000 : _zz_shift_q_0_14 = shift_q_map_24;
      6'b011001 : _zz_shift_q_0_14 = shift_q_map_25;
      6'b011010 : _zz_shift_q_0_14 = shift_q_map_26;
      6'b011011 : _zz_shift_q_0_14 = shift_q_map_27;
      6'b011100 : _zz_shift_q_0_14 = shift_q_map_28;
      6'b011101 : _zz_shift_q_0_14 = shift_q_map_29;
      6'b011110 : _zz_shift_q_0_14 = shift_q_map_30;
      6'b011111 : _zz_shift_q_0_14 = shift_q_map_31;
      6'b100000 : _zz_shift_q_0_14 = shift_q_map_32;
      6'b100001 : _zz_shift_q_0_14 = shift_q_map_33;
      6'b100010 : _zz_shift_q_0_14 = shift_q_map_34;
      6'b100011 : _zz_shift_q_0_14 = shift_q_map_35;
      6'b100100 : _zz_shift_q_0_14 = shift_q_map_36;
      6'b100101 : _zz_shift_q_0_14 = shift_q_map_37;
      6'b100110 : _zz_shift_q_0_14 = shift_q_map_38;
      6'b100111 : _zz_shift_q_0_14 = shift_q_map_39;
      6'b101000 : _zz_shift_q_0_14 = shift_q_map_40;
      6'b101001 : _zz_shift_q_0_14 = shift_q_map_41;
      6'b101010 : _zz_shift_q_0_14 = shift_q_map_42;
      6'b101011 : _zz_shift_q_0_14 = shift_q_map_43;
      6'b101100 : _zz_shift_q_0_14 = shift_q_map_44;
      6'b101101 : _zz_shift_q_0_14 = shift_q_map_45;
      6'b101110 : _zz_shift_q_0_14 = shift_q_map_46;
      6'b101111 : _zz_shift_q_0_14 = shift_q_map_47;
      6'b110000 : _zz_shift_q_0_14 = shift_q_map_48;
      6'b110001 : _zz_shift_q_0_14 = shift_q_map_49;
      6'b110010 : _zz_shift_q_0_14 = shift_q_map_50;
      6'b110011 : _zz_shift_q_0_14 = shift_q_map_51;
      6'b110100 : _zz_shift_q_0_14 = shift_q_map_52;
      6'b110101 : _zz_shift_q_0_14 = shift_q_map_53;
      6'b110110 : _zz_shift_q_0_14 = shift_q_map_54;
      6'b110111 : _zz_shift_q_0_14 = shift_q_map_55;
      6'b111000 : _zz_shift_q_0_14 = shift_q_map_56;
      6'b111001 : _zz_shift_q_0_14 = shift_q_map_57;
      6'b111010 : _zz_shift_q_0_14 = shift_q_map_58;
      6'b111011 : _zz_shift_q_0_14 = shift_q_map_59;
      6'b111100 : _zz_shift_q_0_14 = shift_q_map_60;
      6'b111101 : _zz_shift_q_0_14 = shift_q_map_61;
      6'b111110 : _zz_shift_q_0_14 = shift_q_map_62;
      default : _zz_shift_q_0_14 = shift_q_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_1_15)
      6'b000000 : _zz_shift_i_1_14 = shift_i_map_0;
      6'b000001 : _zz_shift_i_1_14 = shift_i_map_1;
      6'b000010 : _zz_shift_i_1_14 = shift_i_map_2;
      6'b000011 : _zz_shift_i_1_14 = shift_i_map_3;
      6'b000100 : _zz_shift_i_1_14 = shift_i_map_4;
      6'b000101 : _zz_shift_i_1_14 = shift_i_map_5;
      6'b000110 : _zz_shift_i_1_14 = shift_i_map_6;
      6'b000111 : _zz_shift_i_1_14 = shift_i_map_7;
      6'b001000 : _zz_shift_i_1_14 = shift_i_map_8;
      6'b001001 : _zz_shift_i_1_14 = shift_i_map_9;
      6'b001010 : _zz_shift_i_1_14 = shift_i_map_10;
      6'b001011 : _zz_shift_i_1_14 = shift_i_map_11;
      6'b001100 : _zz_shift_i_1_14 = shift_i_map_12;
      6'b001101 : _zz_shift_i_1_14 = shift_i_map_13;
      6'b001110 : _zz_shift_i_1_14 = shift_i_map_14;
      6'b001111 : _zz_shift_i_1_14 = shift_i_map_15;
      6'b010000 : _zz_shift_i_1_14 = shift_i_map_16;
      6'b010001 : _zz_shift_i_1_14 = shift_i_map_17;
      6'b010010 : _zz_shift_i_1_14 = shift_i_map_18;
      6'b010011 : _zz_shift_i_1_14 = shift_i_map_19;
      6'b010100 : _zz_shift_i_1_14 = shift_i_map_20;
      6'b010101 : _zz_shift_i_1_14 = shift_i_map_21;
      6'b010110 : _zz_shift_i_1_14 = shift_i_map_22;
      6'b010111 : _zz_shift_i_1_14 = shift_i_map_23;
      6'b011000 : _zz_shift_i_1_14 = shift_i_map_24;
      6'b011001 : _zz_shift_i_1_14 = shift_i_map_25;
      6'b011010 : _zz_shift_i_1_14 = shift_i_map_26;
      6'b011011 : _zz_shift_i_1_14 = shift_i_map_27;
      6'b011100 : _zz_shift_i_1_14 = shift_i_map_28;
      6'b011101 : _zz_shift_i_1_14 = shift_i_map_29;
      6'b011110 : _zz_shift_i_1_14 = shift_i_map_30;
      6'b011111 : _zz_shift_i_1_14 = shift_i_map_31;
      6'b100000 : _zz_shift_i_1_14 = shift_i_map_32;
      6'b100001 : _zz_shift_i_1_14 = shift_i_map_33;
      6'b100010 : _zz_shift_i_1_14 = shift_i_map_34;
      6'b100011 : _zz_shift_i_1_14 = shift_i_map_35;
      6'b100100 : _zz_shift_i_1_14 = shift_i_map_36;
      6'b100101 : _zz_shift_i_1_14 = shift_i_map_37;
      6'b100110 : _zz_shift_i_1_14 = shift_i_map_38;
      6'b100111 : _zz_shift_i_1_14 = shift_i_map_39;
      6'b101000 : _zz_shift_i_1_14 = shift_i_map_40;
      6'b101001 : _zz_shift_i_1_14 = shift_i_map_41;
      6'b101010 : _zz_shift_i_1_14 = shift_i_map_42;
      6'b101011 : _zz_shift_i_1_14 = shift_i_map_43;
      6'b101100 : _zz_shift_i_1_14 = shift_i_map_44;
      6'b101101 : _zz_shift_i_1_14 = shift_i_map_45;
      6'b101110 : _zz_shift_i_1_14 = shift_i_map_46;
      6'b101111 : _zz_shift_i_1_14 = shift_i_map_47;
      6'b110000 : _zz_shift_i_1_14 = shift_i_map_48;
      6'b110001 : _zz_shift_i_1_14 = shift_i_map_49;
      6'b110010 : _zz_shift_i_1_14 = shift_i_map_50;
      6'b110011 : _zz_shift_i_1_14 = shift_i_map_51;
      6'b110100 : _zz_shift_i_1_14 = shift_i_map_52;
      6'b110101 : _zz_shift_i_1_14 = shift_i_map_53;
      6'b110110 : _zz_shift_i_1_14 = shift_i_map_54;
      6'b110111 : _zz_shift_i_1_14 = shift_i_map_55;
      6'b111000 : _zz_shift_i_1_14 = shift_i_map_56;
      6'b111001 : _zz_shift_i_1_14 = shift_i_map_57;
      6'b111010 : _zz_shift_i_1_14 = shift_i_map_58;
      6'b111011 : _zz_shift_i_1_14 = shift_i_map_59;
      6'b111100 : _zz_shift_i_1_14 = shift_i_map_60;
      6'b111101 : _zz_shift_i_1_14 = shift_i_map_61;
      6'b111110 : _zz_shift_i_1_14 = shift_i_map_62;
      default : _zz_shift_i_1_14 = shift_i_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_1_15)
      6'b000000 : _zz_shift_q_1_14 = shift_q_map_0;
      6'b000001 : _zz_shift_q_1_14 = shift_q_map_1;
      6'b000010 : _zz_shift_q_1_14 = shift_q_map_2;
      6'b000011 : _zz_shift_q_1_14 = shift_q_map_3;
      6'b000100 : _zz_shift_q_1_14 = shift_q_map_4;
      6'b000101 : _zz_shift_q_1_14 = shift_q_map_5;
      6'b000110 : _zz_shift_q_1_14 = shift_q_map_6;
      6'b000111 : _zz_shift_q_1_14 = shift_q_map_7;
      6'b001000 : _zz_shift_q_1_14 = shift_q_map_8;
      6'b001001 : _zz_shift_q_1_14 = shift_q_map_9;
      6'b001010 : _zz_shift_q_1_14 = shift_q_map_10;
      6'b001011 : _zz_shift_q_1_14 = shift_q_map_11;
      6'b001100 : _zz_shift_q_1_14 = shift_q_map_12;
      6'b001101 : _zz_shift_q_1_14 = shift_q_map_13;
      6'b001110 : _zz_shift_q_1_14 = shift_q_map_14;
      6'b001111 : _zz_shift_q_1_14 = shift_q_map_15;
      6'b010000 : _zz_shift_q_1_14 = shift_q_map_16;
      6'b010001 : _zz_shift_q_1_14 = shift_q_map_17;
      6'b010010 : _zz_shift_q_1_14 = shift_q_map_18;
      6'b010011 : _zz_shift_q_1_14 = shift_q_map_19;
      6'b010100 : _zz_shift_q_1_14 = shift_q_map_20;
      6'b010101 : _zz_shift_q_1_14 = shift_q_map_21;
      6'b010110 : _zz_shift_q_1_14 = shift_q_map_22;
      6'b010111 : _zz_shift_q_1_14 = shift_q_map_23;
      6'b011000 : _zz_shift_q_1_14 = shift_q_map_24;
      6'b011001 : _zz_shift_q_1_14 = shift_q_map_25;
      6'b011010 : _zz_shift_q_1_14 = shift_q_map_26;
      6'b011011 : _zz_shift_q_1_14 = shift_q_map_27;
      6'b011100 : _zz_shift_q_1_14 = shift_q_map_28;
      6'b011101 : _zz_shift_q_1_14 = shift_q_map_29;
      6'b011110 : _zz_shift_q_1_14 = shift_q_map_30;
      6'b011111 : _zz_shift_q_1_14 = shift_q_map_31;
      6'b100000 : _zz_shift_q_1_14 = shift_q_map_32;
      6'b100001 : _zz_shift_q_1_14 = shift_q_map_33;
      6'b100010 : _zz_shift_q_1_14 = shift_q_map_34;
      6'b100011 : _zz_shift_q_1_14 = shift_q_map_35;
      6'b100100 : _zz_shift_q_1_14 = shift_q_map_36;
      6'b100101 : _zz_shift_q_1_14 = shift_q_map_37;
      6'b100110 : _zz_shift_q_1_14 = shift_q_map_38;
      6'b100111 : _zz_shift_q_1_14 = shift_q_map_39;
      6'b101000 : _zz_shift_q_1_14 = shift_q_map_40;
      6'b101001 : _zz_shift_q_1_14 = shift_q_map_41;
      6'b101010 : _zz_shift_q_1_14 = shift_q_map_42;
      6'b101011 : _zz_shift_q_1_14 = shift_q_map_43;
      6'b101100 : _zz_shift_q_1_14 = shift_q_map_44;
      6'b101101 : _zz_shift_q_1_14 = shift_q_map_45;
      6'b101110 : _zz_shift_q_1_14 = shift_q_map_46;
      6'b101111 : _zz_shift_q_1_14 = shift_q_map_47;
      6'b110000 : _zz_shift_q_1_14 = shift_q_map_48;
      6'b110001 : _zz_shift_q_1_14 = shift_q_map_49;
      6'b110010 : _zz_shift_q_1_14 = shift_q_map_50;
      6'b110011 : _zz_shift_q_1_14 = shift_q_map_51;
      6'b110100 : _zz_shift_q_1_14 = shift_q_map_52;
      6'b110101 : _zz_shift_q_1_14 = shift_q_map_53;
      6'b110110 : _zz_shift_q_1_14 = shift_q_map_54;
      6'b110111 : _zz_shift_q_1_14 = shift_q_map_55;
      6'b111000 : _zz_shift_q_1_14 = shift_q_map_56;
      6'b111001 : _zz_shift_q_1_14 = shift_q_map_57;
      6'b111010 : _zz_shift_q_1_14 = shift_q_map_58;
      6'b111011 : _zz_shift_q_1_14 = shift_q_map_59;
      6'b111100 : _zz_shift_q_1_14 = shift_q_map_60;
      6'b111101 : _zz_shift_q_1_14 = shift_q_map_61;
      6'b111110 : _zz_shift_q_1_14 = shift_q_map_62;
      default : _zz_shift_q_1_14 = shift_q_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_2_15)
      6'b000000 : _zz_shift_i_2_14 = shift_i_map_0;
      6'b000001 : _zz_shift_i_2_14 = shift_i_map_1;
      6'b000010 : _zz_shift_i_2_14 = shift_i_map_2;
      6'b000011 : _zz_shift_i_2_14 = shift_i_map_3;
      6'b000100 : _zz_shift_i_2_14 = shift_i_map_4;
      6'b000101 : _zz_shift_i_2_14 = shift_i_map_5;
      6'b000110 : _zz_shift_i_2_14 = shift_i_map_6;
      6'b000111 : _zz_shift_i_2_14 = shift_i_map_7;
      6'b001000 : _zz_shift_i_2_14 = shift_i_map_8;
      6'b001001 : _zz_shift_i_2_14 = shift_i_map_9;
      6'b001010 : _zz_shift_i_2_14 = shift_i_map_10;
      6'b001011 : _zz_shift_i_2_14 = shift_i_map_11;
      6'b001100 : _zz_shift_i_2_14 = shift_i_map_12;
      6'b001101 : _zz_shift_i_2_14 = shift_i_map_13;
      6'b001110 : _zz_shift_i_2_14 = shift_i_map_14;
      6'b001111 : _zz_shift_i_2_14 = shift_i_map_15;
      6'b010000 : _zz_shift_i_2_14 = shift_i_map_16;
      6'b010001 : _zz_shift_i_2_14 = shift_i_map_17;
      6'b010010 : _zz_shift_i_2_14 = shift_i_map_18;
      6'b010011 : _zz_shift_i_2_14 = shift_i_map_19;
      6'b010100 : _zz_shift_i_2_14 = shift_i_map_20;
      6'b010101 : _zz_shift_i_2_14 = shift_i_map_21;
      6'b010110 : _zz_shift_i_2_14 = shift_i_map_22;
      6'b010111 : _zz_shift_i_2_14 = shift_i_map_23;
      6'b011000 : _zz_shift_i_2_14 = shift_i_map_24;
      6'b011001 : _zz_shift_i_2_14 = shift_i_map_25;
      6'b011010 : _zz_shift_i_2_14 = shift_i_map_26;
      6'b011011 : _zz_shift_i_2_14 = shift_i_map_27;
      6'b011100 : _zz_shift_i_2_14 = shift_i_map_28;
      6'b011101 : _zz_shift_i_2_14 = shift_i_map_29;
      6'b011110 : _zz_shift_i_2_14 = shift_i_map_30;
      6'b011111 : _zz_shift_i_2_14 = shift_i_map_31;
      6'b100000 : _zz_shift_i_2_14 = shift_i_map_32;
      6'b100001 : _zz_shift_i_2_14 = shift_i_map_33;
      6'b100010 : _zz_shift_i_2_14 = shift_i_map_34;
      6'b100011 : _zz_shift_i_2_14 = shift_i_map_35;
      6'b100100 : _zz_shift_i_2_14 = shift_i_map_36;
      6'b100101 : _zz_shift_i_2_14 = shift_i_map_37;
      6'b100110 : _zz_shift_i_2_14 = shift_i_map_38;
      6'b100111 : _zz_shift_i_2_14 = shift_i_map_39;
      6'b101000 : _zz_shift_i_2_14 = shift_i_map_40;
      6'b101001 : _zz_shift_i_2_14 = shift_i_map_41;
      6'b101010 : _zz_shift_i_2_14 = shift_i_map_42;
      6'b101011 : _zz_shift_i_2_14 = shift_i_map_43;
      6'b101100 : _zz_shift_i_2_14 = shift_i_map_44;
      6'b101101 : _zz_shift_i_2_14 = shift_i_map_45;
      6'b101110 : _zz_shift_i_2_14 = shift_i_map_46;
      6'b101111 : _zz_shift_i_2_14 = shift_i_map_47;
      6'b110000 : _zz_shift_i_2_14 = shift_i_map_48;
      6'b110001 : _zz_shift_i_2_14 = shift_i_map_49;
      6'b110010 : _zz_shift_i_2_14 = shift_i_map_50;
      6'b110011 : _zz_shift_i_2_14 = shift_i_map_51;
      6'b110100 : _zz_shift_i_2_14 = shift_i_map_52;
      6'b110101 : _zz_shift_i_2_14 = shift_i_map_53;
      6'b110110 : _zz_shift_i_2_14 = shift_i_map_54;
      6'b110111 : _zz_shift_i_2_14 = shift_i_map_55;
      6'b111000 : _zz_shift_i_2_14 = shift_i_map_56;
      6'b111001 : _zz_shift_i_2_14 = shift_i_map_57;
      6'b111010 : _zz_shift_i_2_14 = shift_i_map_58;
      6'b111011 : _zz_shift_i_2_14 = shift_i_map_59;
      6'b111100 : _zz_shift_i_2_14 = shift_i_map_60;
      6'b111101 : _zz_shift_i_2_14 = shift_i_map_61;
      6'b111110 : _zz_shift_i_2_14 = shift_i_map_62;
      default : _zz_shift_i_2_14 = shift_i_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_2_15)
      6'b000000 : _zz_shift_q_2_14 = shift_q_map_0;
      6'b000001 : _zz_shift_q_2_14 = shift_q_map_1;
      6'b000010 : _zz_shift_q_2_14 = shift_q_map_2;
      6'b000011 : _zz_shift_q_2_14 = shift_q_map_3;
      6'b000100 : _zz_shift_q_2_14 = shift_q_map_4;
      6'b000101 : _zz_shift_q_2_14 = shift_q_map_5;
      6'b000110 : _zz_shift_q_2_14 = shift_q_map_6;
      6'b000111 : _zz_shift_q_2_14 = shift_q_map_7;
      6'b001000 : _zz_shift_q_2_14 = shift_q_map_8;
      6'b001001 : _zz_shift_q_2_14 = shift_q_map_9;
      6'b001010 : _zz_shift_q_2_14 = shift_q_map_10;
      6'b001011 : _zz_shift_q_2_14 = shift_q_map_11;
      6'b001100 : _zz_shift_q_2_14 = shift_q_map_12;
      6'b001101 : _zz_shift_q_2_14 = shift_q_map_13;
      6'b001110 : _zz_shift_q_2_14 = shift_q_map_14;
      6'b001111 : _zz_shift_q_2_14 = shift_q_map_15;
      6'b010000 : _zz_shift_q_2_14 = shift_q_map_16;
      6'b010001 : _zz_shift_q_2_14 = shift_q_map_17;
      6'b010010 : _zz_shift_q_2_14 = shift_q_map_18;
      6'b010011 : _zz_shift_q_2_14 = shift_q_map_19;
      6'b010100 : _zz_shift_q_2_14 = shift_q_map_20;
      6'b010101 : _zz_shift_q_2_14 = shift_q_map_21;
      6'b010110 : _zz_shift_q_2_14 = shift_q_map_22;
      6'b010111 : _zz_shift_q_2_14 = shift_q_map_23;
      6'b011000 : _zz_shift_q_2_14 = shift_q_map_24;
      6'b011001 : _zz_shift_q_2_14 = shift_q_map_25;
      6'b011010 : _zz_shift_q_2_14 = shift_q_map_26;
      6'b011011 : _zz_shift_q_2_14 = shift_q_map_27;
      6'b011100 : _zz_shift_q_2_14 = shift_q_map_28;
      6'b011101 : _zz_shift_q_2_14 = shift_q_map_29;
      6'b011110 : _zz_shift_q_2_14 = shift_q_map_30;
      6'b011111 : _zz_shift_q_2_14 = shift_q_map_31;
      6'b100000 : _zz_shift_q_2_14 = shift_q_map_32;
      6'b100001 : _zz_shift_q_2_14 = shift_q_map_33;
      6'b100010 : _zz_shift_q_2_14 = shift_q_map_34;
      6'b100011 : _zz_shift_q_2_14 = shift_q_map_35;
      6'b100100 : _zz_shift_q_2_14 = shift_q_map_36;
      6'b100101 : _zz_shift_q_2_14 = shift_q_map_37;
      6'b100110 : _zz_shift_q_2_14 = shift_q_map_38;
      6'b100111 : _zz_shift_q_2_14 = shift_q_map_39;
      6'b101000 : _zz_shift_q_2_14 = shift_q_map_40;
      6'b101001 : _zz_shift_q_2_14 = shift_q_map_41;
      6'b101010 : _zz_shift_q_2_14 = shift_q_map_42;
      6'b101011 : _zz_shift_q_2_14 = shift_q_map_43;
      6'b101100 : _zz_shift_q_2_14 = shift_q_map_44;
      6'b101101 : _zz_shift_q_2_14 = shift_q_map_45;
      6'b101110 : _zz_shift_q_2_14 = shift_q_map_46;
      6'b101111 : _zz_shift_q_2_14 = shift_q_map_47;
      6'b110000 : _zz_shift_q_2_14 = shift_q_map_48;
      6'b110001 : _zz_shift_q_2_14 = shift_q_map_49;
      6'b110010 : _zz_shift_q_2_14 = shift_q_map_50;
      6'b110011 : _zz_shift_q_2_14 = shift_q_map_51;
      6'b110100 : _zz_shift_q_2_14 = shift_q_map_52;
      6'b110101 : _zz_shift_q_2_14 = shift_q_map_53;
      6'b110110 : _zz_shift_q_2_14 = shift_q_map_54;
      6'b110111 : _zz_shift_q_2_14 = shift_q_map_55;
      6'b111000 : _zz_shift_q_2_14 = shift_q_map_56;
      6'b111001 : _zz_shift_q_2_14 = shift_q_map_57;
      6'b111010 : _zz_shift_q_2_14 = shift_q_map_58;
      6'b111011 : _zz_shift_q_2_14 = shift_q_map_59;
      6'b111100 : _zz_shift_q_2_14 = shift_q_map_60;
      6'b111101 : _zz_shift_q_2_14 = shift_q_map_61;
      6'b111110 : _zz_shift_q_2_14 = shift_q_map_62;
      default : _zz_shift_q_2_14 = shift_q_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_3_15)
      6'b000000 : _zz_shift_i_3_14 = shift_i_map_0;
      6'b000001 : _zz_shift_i_3_14 = shift_i_map_1;
      6'b000010 : _zz_shift_i_3_14 = shift_i_map_2;
      6'b000011 : _zz_shift_i_3_14 = shift_i_map_3;
      6'b000100 : _zz_shift_i_3_14 = shift_i_map_4;
      6'b000101 : _zz_shift_i_3_14 = shift_i_map_5;
      6'b000110 : _zz_shift_i_3_14 = shift_i_map_6;
      6'b000111 : _zz_shift_i_3_14 = shift_i_map_7;
      6'b001000 : _zz_shift_i_3_14 = shift_i_map_8;
      6'b001001 : _zz_shift_i_3_14 = shift_i_map_9;
      6'b001010 : _zz_shift_i_3_14 = shift_i_map_10;
      6'b001011 : _zz_shift_i_3_14 = shift_i_map_11;
      6'b001100 : _zz_shift_i_3_14 = shift_i_map_12;
      6'b001101 : _zz_shift_i_3_14 = shift_i_map_13;
      6'b001110 : _zz_shift_i_3_14 = shift_i_map_14;
      6'b001111 : _zz_shift_i_3_14 = shift_i_map_15;
      6'b010000 : _zz_shift_i_3_14 = shift_i_map_16;
      6'b010001 : _zz_shift_i_3_14 = shift_i_map_17;
      6'b010010 : _zz_shift_i_3_14 = shift_i_map_18;
      6'b010011 : _zz_shift_i_3_14 = shift_i_map_19;
      6'b010100 : _zz_shift_i_3_14 = shift_i_map_20;
      6'b010101 : _zz_shift_i_3_14 = shift_i_map_21;
      6'b010110 : _zz_shift_i_3_14 = shift_i_map_22;
      6'b010111 : _zz_shift_i_3_14 = shift_i_map_23;
      6'b011000 : _zz_shift_i_3_14 = shift_i_map_24;
      6'b011001 : _zz_shift_i_3_14 = shift_i_map_25;
      6'b011010 : _zz_shift_i_3_14 = shift_i_map_26;
      6'b011011 : _zz_shift_i_3_14 = shift_i_map_27;
      6'b011100 : _zz_shift_i_3_14 = shift_i_map_28;
      6'b011101 : _zz_shift_i_3_14 = shift_i_map_29;
      6'b011110 : _zz_shift_i_3_14 = shift_i_map_30;
      6'b011111 : _zz_shift_i_3_14 = shift_i_map_31;
      6'b100000 : _zz_shift_i_3_14 = shift_i_map_32;
      6'b100001 : _zz_shift_i_3_14 = shift_i_map_33;
      6'b100010 : _zz_shift_i_3_14 = shift_i_map_34;
      6'b100011 : _zz_shift_i_3_14 = shift_i_map_35;
      6'b100100 : _zz_shift_i_3_14 = shift_i_map_36;
      6'b100101 : _zz_shift_i_3_14 = shift_i_map_37;
      6'b100110 : _zz_shift_i_3_14 = shift_i_map_38;
      6'b100111 : _zz_shift_i_3_14 = shift_i_map_39;
      6'b101000 : _zz_shift_i_3_14 = shift_i_map_40;
      6'b101001 : _zz_shift_i_3_14 = shift_i_map_41;
      6'b101010 : _zz_shift_i_3_14 = shift_i_map_42;
      6'b101011 : _zz_shift_i_3_14 = shift_i_map_43;
      6'b101100 : _zz_shift_i_3_14 = shift_i_map_44;
      6'b101101 : _zz_shift_i_3_14 = shift_i_map_45;
      6'b101110 : _zz_shift_i_3_14 = shift_i_map_46;
      6'b101111 : _zz_shift_i_3_14 = shift_i_map_47;
      6'b110000 : _zz_shift_i_3_14 = shift_i_map_48;
      6'b110001 : _zz_shift_i_3_14 = shift_i_map_49;
      6'b110010 : _zz_shift_i_3_14 = shift_i_map_50;
      6'b110011 : _zz_shift_i_3_14 = shift_i_map_51;
      6'b110100 : _zz_shift_i_3_14 = shift_i_map_52;
      6'b110101 : _zz_shift_i_3_14 = shift_i_map_53;
      6'b110110 : _zz_shift_i_3_14 = shift_i_map_54;
      6'b110111 : _zz_shift_i_3_14 = shift_i_map_55;
      6'b111000 : _zz_shift_i_3_14 = shift_i_map_56;
      6'b111001 : _zz_shift_i_3_14 = shift_i_map_57;
      6'b111010 : _zz_shift_i_3_14 = shift_i_map_58;
      6'b111011 : _zz_shift_i_3_14 = shift_i_map_59;
      6'b111100 : _zz_shift_i_3_14 = shift_i_map_60;
      6'b111101 : _zz_shift_i_3_14 = shift_i_map_61;
      6'b111110 : _zz_shift_i_3_14 = shift_i_map_62;
      default : _zz_shift_i_3_14 = shift_i_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_3_15)
      6'b000000 : _zz_shift_q_3_14 = shift_q_map_0;
      6'b000001 : _zz_shift_q_3_14 = shift_q_map_1;
      6'b000010 : _zz_shift_q_3_14 = shift_q_map_2;
      6'b000011 : _zz_shift_q_3_14 = shift_q_map_3;
      6'b000100 : _zz_shift_q_3_14 = shift_q_map_4;
      6'b000101 : _zz_shift_q_3_14 = shift_q_map_5;
      6'b000110 : _zz_shift_q_3_14 = shift_q_map_6;
      6'b000111 : _zz_shift_q_3_14 = shift_q_map_7;
      6'b001000 : _zz_shift_q_3_14 = shift_q_map_8;
      6'b001001 : _zz_shift_q_3_14 = shift_q_map_9;
      6'b001010 : _zz_shift_q_3_14 = shift_q_map_10;
      6'b001011 : _zz_shift_q_3_14 = shift_q_map_11;
      6'b001100 : _zz_shift_q_3_14 = shift_q_map_12;
      6'b001101 : _zz_shift_q_3_14 = shift_q_map_13;
      6'b001110 : _zz_shift_q_3_14 = shift_q_map_14;
      6'b001111 : _zz_shift_q_3_14 = shift_q_map_15;
      6'b010000 : _zz_shift_q_3_14 = shift_q_map_16;
      6'b010001 : _zz_shift_q_3_14 = shift_q_map_17;
      6'b010010 : _zz_shift_q_3_14 = shift_q_map_18;
      6'b010011 : _zz_shift_q_3_14 = shift_q_map_19;
      6'b010100 : _zz_shift_q_3_14 = shift_q_map_20;
      6'b010101 : _zz_shift_q_3_14 = shift_q_map_21;
      6'b010110 : _zz_shift_q_3_14 = shift_q_map_22;
      6'b010111 : _zz_shift_q_3_14 = shift_q_map_23;
      6'b011000 : _zz_shift_q_3_14 = shift_q_map_24;
      6'b011001 : _zz_shift_q_3_14 = shift_q_map_25;
      6'b011010 : _zz_shift_q_3_14 = shift_q_map_26;
      6'b011011 : _zz_shift_q_3_14 = shift_q_map_27;
      6'b011100 : _zz_shift_q_3_14 = shift_q_map_28;
      6'b011101 : _zz_shift_q_3_14 = shift_q_map_29;
      6'b011110 : _zz_shift_q_3_14 = shift_q_map_30;
      6'b011111 : _zz_shift_q_3_14 = shift_q_map_31;
      6'b100000 : _zz_shift_q_3_14 = shift_q_map_32;
      6'b100001 : _zz_shift_q_3_14 = shift_q_map_33;
      6'b100010 : _zz_shift_q_3_14 = shift_q_map_34;
      6'b100011 : _zz_shift_q_3_14 = shift_q_map_35;
      6'b100100 : _zz_shift_q_3_14 = shift_q_map_36;
      6'b100101 : _zz_shift_q_3_14 = shift_q_map_37;
      6'b100110 : _zz_shift_q_3_14 = shift_q_map_38;
      6'b100111 : _zz_shift_q_3_14 = shift_q_map_39;
      6'b101000 : _zz_shift_q_3_14 = shift_q_map_40;
      6'b101001 : _zz_shift_q_3_14 = shift_q_map_41;
      6'b101010 : _zz_shift_q_3_14 = shift_q_map_42;
      6'b101011 : _zz_shift_q_3_14 = shift_q_map_43;
      6'b101100 : _zz_shift_q_3_14 = shift_q_map_44;
      6'b101101 : _zz_shift_q_3_14 = shift_q_map_45;
      6'b101110 : _zz_shift_q_3_14 = shift_q_map_46;
      6'b101111 : _zz_shift_q_3_14 = shift_q_map_47;
      6'b110000 : _zz_shift_q_3_14 = shift_q_map_48;
      6'b110001 : _zz_shift_q_3_14 = shift_q_map_49;
      6'b110010 : _zz_shift_q_3_14 = shift_q_map_50;
      6'b110011 : _zz_shift_q_3_14 = shift_q_map_51;
      6'b110100 : _zz_shift_q_3_14 = shift_q_map_52;
      6'b110101 : _zz_shift_q_3_14 = shift_q_map_53;
      6'b110110 : _zz_shift_q_3_14 = shift_q_map_54;
      6'b110111 : _zz_shift_q_3_14 = shift_q_map_55;
      6'b111000 : _zz_shift_q_3_14 = shift_q_map_56;
      6'b111001 : _zz_shift_q_3_14 = shift_q_map_57;
      6'b111010 : _zz_shift_q_3_14 = shift_q_map_58;
      6'b111011 : _zz_shift_q_3_14 = shift_q_map_59;
      6'b111100 : _zz_shift_q_3_14 = shift_q_map_60;
      6'b111101 : _zz_shift_q_3_14 = shift_q_map_61;
      6'b111110 : _zz_shift_q_3_14 = shift_q_map_62;
      default : _zz_shift_q_3_14 = shift_q_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_4_15)
      6'b000000 : _zz_shift_i_4_14 = shift_i_map_0;
      6'b000001 : _zz_shift_i_4_14 = shift_i_map_1;
      6'b000010 : _zz_shift_i_4_14 = shift_i_map_2;
      6'b000011 : _zz_shift_i_4_14 = shift_i_map_3;
      6'b000100 : _zz_shift_i_4_14 = shift_i_map_4;
      6'b000101 : _zz_shift_i_4_14 = shift_i_map_5;
      6'b000110 : _zz_shift_i_4_14 = shift_i_map_6;
      6'b000111 : _zz_shift_i_4_14 = shift_i_map_7;
      6'b001000 : _zz_shift_i_4_14 = shift_i_map_8;
      6'b001001 : _zz_shift_i_4_14 = shift_i_map_9;
      6'b001010 : _zz_shift_i_4_14 = shift_i_map_10;
      6'b001011 : _zz_shift_i_4_14 = shift_i_map_11;
      6'b001100 : _zz_shift_i_4_14 = shift_i_map_12;
      6'b001101 : _zz_shift_i_4_14 = shift_i_map_13;
      6'b001110 : _zz_shift_i_4_14 = shift_i_map_14;
      6'b001111 : _zz_shift_i_4_14 = shift_i_map_15;
      6'b010000 : _zz_shift_i_4_14 = shift_i_map_16;
      6'b010001 : _zz_shift_i_4_14 = shift_i_map_17;
      6'b010010 : _zz_shift_i_4_14 = shift_i_map_18;
      6'b010011 : _zz_shift_i_4_14 = shift_i_map_19;
      6'b010100 : _zz_shift_i_4_14 = shift_i_map_20;
      6'b010101 : _zz_shift_i_4_14 = shift_i_map_21;
      6'b010110 : _zz_shift_i_4_14 = shift_i_map_22;
      6'b010111 : _zz_shift_i_4_14 = shift_i_map_23;
      6'b011000 : _zz_shift_i_4_14 = shift_i_map_24;
      6'b011001 : _zz_shift_i_4_14 = shift_i_map_25;
      6'b011010 : _zz_shift_i_4_14 = shift_i_map_26;
      6'b011011 : _zz_shift_i_4_14 = shift_i_map_27;
      6'b011100 : _zz_shift_i_4_14 = shift_i_map_28;
      6'b011101 : _zz_shift_i_4_14 = shift_i_map_29;
      6'b011110 : _zz_shift_i_4_14 = shift_i_map_30;
      6'b011111 : _zz_shift_i_4_14 = shift_i_map_31;
      6'b100000 : _zz_shift_i_4_14 = shift_i_map_32;
      6'b100001 : _zz_shift_i_4_14 = shift_i_map_33;
      6'b100010 : _zz_shift_i_4_14 = shift_i_map_34;
      6'b100011 : _zz_shift_i_4_14 = shift_i_map_35;
      6'b100100 : _zz_shift_i_4_14 = shift_i_map_36;
      6'b100101 : _zz_shift_i_4_14 = shift_i_map_37;
      6'b100110 : _zz_shift_i_4_14 = shift_i_map_38;
      6'b100111 : _zz_shift_i_4_14 = shift_i_map_39;
      6'b101000 : _zz_shift_i_4_14 = shift_i_map_40;
      6'b101001 : _zz_shift_i_4_14 = shift_i_map_41;
      6'b101010 : _zz_shift_i_4_14 = shift_i_map_42;
      6'b101011 : _zz_shift_i_4_14 = shift_i_map_43;
      6'b101100 : _zz_shift_i_4_14 = shift_i_map_44;
      6'b101101 : _zz_shift_i_4_14 = shift_i_map_45;
      6'b101110 : _zz_shift_i_4_14 = shift_i_map_46;
      6'b101111 : _zz_shift_i_4_14 = shift_i_map_47;
      6'b110000 : _zz_shift_i_4_14 = shift_i_map_48;
      6'b110001 : _zz_shift_i_4_14 = shift_i_map_49;
      6'b110010 : _zz_shift_i_4_14 = shift_i_map_50;
      6'b110011 : _zz_shift_i_4_14 = shift_i_map_51;
      6'b110100 : _zz_shift_i_4_14 = shift_i_map_52;
      6'b110101 : _zz_shift_i_4_14 = shift_i_map_53;
      6'b110110 : _zz_shift_i_4_14 = shift_i_map_54;
      6'b110111 : _zz_shift_i_4_14 = shift_i_map_55;
      6'b111000 : _zz_shift_i_4_14 = shift_i_map_56;
      6'b111001 : _zz_shift_i_4_14 = shift_i_map_57;
      6'b111010 : _zz_shift_i_4_14 = shift_i_map_58;
      6'b111011 : _zz_shift_i_4_14 = shift_i_map_59;
      6'b111100 : _zz_shift_i_4_14 = shift_i_map_60;
      6'b111101 : _zz_shift_i_4_14 = shift_i_map_61;
      6'b111110 : _zz_shift_i_4_14 = shift_i_map_62;
      default : _zz_shift_i_4_14 = shift_i_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_4_15)
      6'b000000 : _zz_shift_q_4_14 = shift_q_map_0;
      6'b000001 : _zz_shift_q_4_14 = shift_q_map_1;
      6'b000010 : _zz_shift_q_4_14 = shift_q_map_2;
      6'b000011 : _zz_shift_q_4_14 = shift_q_map_3;
      6'b000100 : _zz_shift_q_4_14 = shift_q_map_4;
      6'b000101 : _zz_shift_q_4_14 = shift_q_map_5;
      6'b000110 : _zz_shift_q_4_14 = shift_q_map_6;
      6'b000111 : _zz_shift_q_4_14 = shift_q_map_7;
      6'b001000 : _zz_shift_q_4_14 = shift_q_map_8;
      6'b001001 : _zz_shift_q_4_14 = shift_q_map_9;
      6'b001010 : _zz_shift_q_4_14 = shift_q_map_10;
      6'b001011 : _zz_shift_q_4_14 = shift_q_map_11;
      6'b001100 : _zz_shift_q_4_14 = shift_q_map_12;
      6'b001101 : _zz_shift_q_4_14 = shift_q_map_13;
      6'b001110 : _zz_shift_q_4_14 = shift_q_map_14;
      6'b001111 : _zz_shift_q_4_14 = shift_q_map_15;
      6'b010000 : _zz_shift_q_4_14 = shift_q_map_16;
      6'b010001 : _zz_shift_q_4_14 = shift_q_map_17;
      6'b010010 : _zz_shift_q_4_14 = shift_q_map_18;
      6'b010011 : _zz_shift_q_4_14 = shift_q_map_19;
      6'b010100 : _zz_shift_q_4_14 = shift_q_map_20;
      6'b010101 : _zz_shift_q_4_14 = shift_q_map_21;
      6'b010110 : _zz_shift_q_4_14 = shift_q_map_22;
      6'b010111 : _zz_shift_q_4_14 = shift_q_map_23;
      6'b011000 : _zz_shift_q_4_14 = shift_q_map_24;
      6'b011001 : _zz_shift_q_4_14 = shift_q_map_25;
      6'b011010 : _zz_shift_q_4_14 = shift_q_map_26;
      6'b011011 : _zz_shift_q_4_14 = shift_q_map_27;
      6'b011100 : _zz_shift_q_4_14 = shift_q_map_28;
      6'b011101 : _zz_shift_q_4_14 = shift_q_map_29;
      6'b011110 : _zz_shift_q_4_14 = shift_q_map_30;
      6'b011111 : _zz_shift_q_4_14 = shift_q_map_31;
      6'b100000 : _zz_shift_q_4_14 = shift_q_map_32;
      6'b100001 : _zz_shift_q_4_14 = shift_q_map_33;
      6'b100010 : _zz_shift_q_4_14 = shift_q_map_34;
      6'b100011 : _zz_shift_q_4_14 = shift_q_map_35;
      6'b100100 : _zz_shift_q_4_14 = shift_q_map_36;
      6'b100101 : _zz_shift_q_4_14 = shift_q_map_37;
      6'b100110 : _zz_shift_q_4_14 = shift_q_map_38;
      6'b100111 : _zz_shift_q_4_14 = shift_q_map_39;
      6'b101000 : _zz_shift_q_4_14 = shift_q_map_40;
      6'b101001 : _zz_shift_q_4_14 = shift_q_map_41;
      6'b101010 : _zz_shift_q_4_14 = shift_q_map_42;
      6'b101011 : _zz_shift_q_4_14 = shift_q_map_43;
      6'b101100 : _zz_shift_q_4_14 = shift_q_map_44;
      6'b101101 : _zz_shift_q_4_14 = shift_q_map_45;
      6'b101110 : _zz_shift_q_4_14 = shift_q_map_46;
      6'b101111 : _zz_shift_q_4_14 = shift_q_map_47;
      6'b110000 : _zz_shift_q_4_14 = shift_q_map_48;
      6'b110001 : _zz_shift_q_4_14 = shift_q_map_49;
      6'b110010 : _zz_shift_q_4_14 = shift_q_map_50;
      6'b110011 : _zz_shift_q_4_14 = shift_q_map_51;
      6'b110100 : _zz_shift_q_4_14 = shift_q_map_52;
      6'b110101 : _zz_shift_q_4_14 = shift_q_map_53;
      6'b110110 : _zz_shift_q_4_14 = shift_q_map_54;
      6'b110111 : _zz_shift_q_4_14 = shift_q_map_55;
      6'b111000 : _zz_shift_q_4_14 = shift_q_map_56;
      6'b111001 : _zz_shift_q_4_14 = shift_q_map_57;
      6'b111010 : _zz_shift_q_4_14 = shift_q_map_58;
      6'b111011 : _zz_shift_q_4_14 = shift_q_map_59;
      6'b111100 : _zz_shift_q_4_14 = shift_q_map_60;
      6'b111101 : _zz_shift_q_4_14 = shift_q_map_61;
      6'b111110 : _zz_shift_q_4_14 = shift_q_map_62;
      default : _zz_shift_q_4_14 = shift_q_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_5_15)
      6'b000000 : _zz_shift_i_5_14 = shift_i_map_0;
      6'b000001 : _zz_shift_i_5_14 = shift_i_map_1;
      6'b000010 : _zz_shift_i_5_14 = shift_i_map_2;
      6'b000011 : _zz_shift_i_5_14 = shift_i_map_3;
      6'b000100 : _zz_shift_i_5_14 = shift_i_map_4;
      6'b000101 : _zz_shift_i_5_14 = shift_i_map_5;
      6'b000110 : _zz_shift_i_5_14 = shift_i_map_6;
      6'b000111 : _zz_shift_i_5_14 = shift_i_map_7;
      6'b001000 : _zz_shift_i_5_14 = shift_i_map_8;
      6'b001001 : _zz_shift_i_5_14 = shift_i_map_9;
      6'b001010 : _zz_shift_i_5_14 = shift_i_map_10;
      6'b001011 : _zz_shift_i_5_14 = shift_i_map_11;
      6'b001100 : _zz_shift_i_5_14 = shift_i_map_12;
      6'b001101 : _zz_shift_i_5_14 = shift_i_map_13;
      6'b001110 : _zz_shift_i_5_14 = shift_i_map_14;
      6'b001111 : _zz_shift_i_5_14 = shift_i_map_15;
      6'b010000 : _zz_shift_i_5_14 = shift_i_map_16;
      6'b010001 : _zz_shift_i_5_14 = shift_i_map_17;
      6'b010010 : _zz_shift_i_5_14 = shift_i_map_18;
      6'b010011 : _zz_shift_i_5_14 = shift_i_map_19;
      6'b010100 : _zz_shift_i_5_14 = shift_i_map_20;
      6'b010101 : _zz_shift_i_5_14 = shift_i_map_21;
      6'b010110 : _zz_shift_i_5_14 = shift_i_map_22;
      6'b010111 : _zz_shift_i_5_14 = shift_i_map_23;
      6'b011000 : _zz_shift_i_5_14 = shift_i_map_24;
      6'b011001 : _zz_shift_i_5_14 = shift_i_map_25;
      6'b011010 : _zz_shift_i_5_14 = shift_i_map_26;
      6'b011011 : _zz_shift_i_5_14 = shift_i_map_27;
      6'b011100 : _zz_shift_i_5_14 = shift_i_map_28;
      6'b011101 : _zz_shift_i_5_14 = shift_i_map_29;
      6'b011110 : _zz_shift_i_5_14 = shift_i_map_30;
      6'b011111 : _zz_shift_i_5_14 = shift_i_map_31;
      6'b100000 : _zz_shift_i_5_14 = shift_i_map_32;
      6'b100001 : _zz_shift_i_5_14 = shift_i_map_33;
      6'b100010 : _zz_shift_i_5_14 = shift_i_map_34;
      6'b100011 : _zz_shift_i_5_14 = shift_i_map_35;
      6'b100100 : _zz_shift_i_5_14 = shift_i_map_36;
      6'b100101 : _zz_shift_i_5_14 = shift_i_map_37;
      6'b100110 : _zz_shift_i_5_14 = shift_i_map_38;
      6'b100111 : _zz_shift_i_5_14 = shift_i_map_39;
      6'b101000 : _zz_shift_i_5_14 = shift_i_map_40;
      6'b101001 : _zz_shift_i_5_14 = shift_i_map_41;
      6'b101010 : _zz_shift_i_5_14 = shift_i_map_42;
      6'b101011 : _zz_shift_i_5_14 = shift_i_map_43;
      6'b101100 : _zz_shift_i_5_14 = shift_i_map_44;
      6'b101101 : _zz_shift_i_5_14 = shift_i_map_45;
      6'b101110 : _zz_shift_i_5_14 = shift_i_map_46;
      6'b101111 : _zz_shift_i_5_14 = shift_i_map_47;
      6'b110000 : _zz_shift_i_5_14 = shift_i_map_48;
      6'b110001 : _zz_shift_i_5_14 = shift_i_map_49;
      6'b110010 : _zz_shift_i_5_14 = shift_i_map_50;
      6'b110011 : _zz_shift_i_5_14 = shift_i_map_51;
      6'b110100 : _zz_shift_i_5_14 = shift_i_map_52;
      6'b110101 : _zz_shift_i_5_14 = shift_i_map_53;
      6'b110110 : _zz_shift_i_5_14 = shift_i_map_54;
      6'b110111 : _zz_shift_i_5_14 = shift_i_map_55;
      6'b111000 : _zz_shift_i_5_14 = shift_i_map_56;
      6'b111001 : _zz_shift_i_5_14 = shift_i_map_57;
      6'b111010 : _zz_shift_i_5_14 = shift_i_map_58;
      6'b111011 : _zz_shift_i_5_14 = shift_i_map_59;
      6'b111100 : _zz_shift_i_5_14 = shift_i_map_60;
      6'b111101 : _zz_shift_i_5_14 = shift_i_map_61;
      6'b111110 : _zz_shift_i_5_14 = shift_i_map_62;
      default : _zz_shift_i_5_14 = shift_i_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_5_15)
      6'b000000 : _zz_shift_q_5_14 = shift_q_map_0;
      6'b000001 : _zz_shift_q_5_14 = shift_q_map_1;
      6'b000010 : _zz_shift_q_5_14 = shift_q_map_2;
      6'b000011 : _zz_shift_q_5_14 = shift_q_map_3;
      6'b000100 : _zz_shift_q_5_14 = shift_q_map_4;
      6'b000101 : _zz_shift_q_5_14 = shift_q_map_5;
      6'b000110 : _zz_shift_q_5_14 = shift_q_map_6;
      6'b000111 : _zz_shift_q_5_14 = shift_q_map_7;
      6'b001000 : _zz_shift_q_5_14 = shift_q_map_8;
      6'b001001 : _zz_shift_q_5_14 = shift_q_map_9;
      6'b001010 : _zz_shift_q_5_14 = shift_q_map_10;
      6'b001011 : _zz_shift_q_5_14 = shift_q_map_11;
      6'b001100 : _zz_shift_q_5_14 = shift_q_map_12;
      6'b001101 : _zz_shift_q_5_14 = shift_q_map_13;
      6'b001110 : _zz_shift_q_5_14 = shift_q_map_14;
      6'b001111 : _zz_shift_q_5_14 = shift_q_map_15;
      6'b010000 : _zz_shift_q_5_14 = shift_q_map_16;
      6'b010001 : _zz_shift_q_5_14 = shift_q_map_17;
      6'b010010 : _zz_shift_q_5_14 = shift_q_map_18;
      6'b010011 : _zz_shift_q_5_14 = shift_q_map_19;
      6'b010100 : _zz_shift_q_5_14 = shift_q_map_20;
      6'b010101 : _zz_shift_q_5_14 = shift_q_map_21;
      6'b010110 : _zz_shift_q_5_14 = shift_q_map_22;
      6'b010111 : _zz_shift_q_5_14 = shift_q_map_23;
      6'b011000 : _zz_shift_q_5_14 = shift_q_map_24;
      6'b011001 : _zz_shift_q_5_14 = shift_q_map_25;
      6'b011010 : _zz_shift_q_5_14 = shift_q_map_26;
      6'b011011 : _zz_shift_q_5_14 = shift_q_map_27;
      6'b011100 : _zz_shift_q_5_14 = shift_q_map_28;
      6'b011101 : _zz_shift_q_5_14 = shift_q_map_29;
      6'b011110 : _zz_shift_q_5_14 = shift_q_map_30;
      6'b011111 : _zz_shift_q_5_14 = shift_q_map_31;
      6'b100000 : _zz_shift_q_5_14 = shift_q_map_32;
      6'b100001 : _zz_shift_q_5_14 = shift_q_map_33;
      6'b100010 : _zz_shift_q_5_14 = shift_q_map_34;
      6'b100011 : _zz_shift_q_5_14 = shift_q_map_35;
      6'b100100 : _zz_shift_q_5_14 = shift_q_map_36;
      6'b100101 : _zz_shift_q_5_14 = shift_q_map_37;
      6'b100110 : _zz_shift_q_5_14 = shift_q_map_38;
      6'b100111 : _zz_shift_q_5_14 = shift_q_map_39;
      6'b101000 : _zz_shift_q_5_14 = shift_q_map_40;
      6'b101001 : _zz_shift_q_5_14 = shift_q_map_41;
      6'b101010 : _zz_shift_q_5_14 = shift_q_map_42;
      6'b101011 : _zz_shift_q_5_14 = shift_q_map_43;
      6'b101100 : _zz_shift_q_5_14 = shift_q_map_44;
      6'b101101 : _zz_shift_q_5_14 = shift_q_map_45;
      6'b101110 : _zz_shift_q_5_14 = shift_q_map_46;
      6'b101111 : _zz_shift_q_5_14 = shift_q_map_47;
      6'b110000 : _zz_shift_q_5_14 = shift_q_map_48;
      6'b110001 : _zz_shift_q_5_14 = shift_q_map_49;
      6'b110010 : _zz_shift_q_5_14 = shift_q_map_50;
      6'b110011 : _zz_shift_q_5_14 = shift_q_map_51;
      6'b110100 : _zz_shift_q_5_14 = shift_q_map_52;
      6'b110101 : _zz_shift_q_5_14 = shift_q_map_53;
      6'b110110 : _zz_shift_q_5_14 = shift_q_map_54;
      6'b110111 : _zz_shift_q_5_14 = shift_q_map_55;
      6'b111000 : _zz_shift_q_5_14 = shift_q_map_56;
      6'b111001 : _zz_shift_q_5_14 = shift_q_map_57;
      6'b111010 : _zz_shift_q_5_14 = shift_q_map_58;
      6'b111011 : _zz_shift_q_5_14 = shift_q_map_59;
      6'b111100 : _zz_shift_q_5_14 = shift_q_map_60;
      6'b111101 : _zz_shift_q_5_14 = shift_q_map_61;
      6'b111110 : _zz_shift_q_5_14 = shift_q_map_62;
      default : _zz_shift_q_5_14 = shift_q_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_6_15)
      6'b000000 : _zz_shift_i_6_14 = shift_i_map_0;
      6'b000001 : _zz_shift_i_6_14 = shift_i_map_1;
      6'b000010 : _zz_shift_i_6_14 = shift_i_map_2;
      6'b000011 : _zz_shift_i_6_14 = shift_i_map_3;
      6'b000100 : _zz_shift_i_6_14 = shift_i_map_4;
      6'b000101 : _zz_shift_i_6_14 = shift_i_map_5;
      6'b000110 : _zz_shift_i_6_14 = shift_i_map_6;
      6'b000111 : _zz_shift_i_6_14 = shift_i_map_7;
      6'b001000 : _zz_shift_i_6_14 = shift_i_map_8;
      6'b001001 : _zz_shift_i_6_14 = shift_i_map_9;
      6'b001010 : _zz_shift_i_6_14 = shift_i_map_10;
      6'b001011 : _zz_shift_i_6_14 = shift_i_map_11;
      6'b001100 : _zz_shift_i_6_14 = shift_i_map_12;
      6'b001101 : _zz_shift_i_6_14 = shift_i_map_13;
      6'b001110 : _zz_shift_i_6_14 = shift_i_map_14;
      6'b001111 : _zz_shift_i_6_14 = shift_i_map_15;
      6'b010000 : _zz_shift_i_6_14 = shift_i_map_16;
      6'b010001 : _zz_shift_i_6_14 = shift_i_map_17;
      6'b010010 : _zz_shift_i_6_14 = shift_i_map_18;
      6'b010011 : _zz_shift_i_6_14 = shift_i_map_19;
      6'b010100 : _zz_shift_i_6_14 = shift_i_map_20;
      6'b010101 : _zz_shift_i_6_14 = shift_i_map_21;
      6'b010110 : _zz_shift_i_6_14 = shift_i_map_22;
      6'b010111 : _zz_shift_i_6_14 = shift_i_map_23;
      6'b011000 : _zz_shift_i_6_14 = shift_i_map_24;
      6'b011001 : _zz_shift_i_6_14 = shift_i_map_25;
      6'b011010 : _zz_shift_i_6_14 = shift_i_map_26;
      6'b011011 : _zz_shift_i_6_14 = shift_i_map_27;
      6'b011100 : _zz_shift_i_6_14 = shift_i_map_28;
      6'b011101 : _zz_shift_i_6_14 = shift_i_map_29;
      6'b011110 : _zz_shift_i_6_14 = shift_i_map_30;
      6'b011111 : _zz_shift_i_6_14 = shift_i_map_31;
      6'b100000 : _zz_shift_i_6_14 = shift_i_map_32;
      6'b100001 : _zz_shift_i_6_14 = shift_i_map_33;
      6'b100010 : _zz_shift_i_6_14 = shift_i_map_34;
      6'b100011 : _zz_shift_i_6_14 = shift_i_map_35;
      6'b100100 : _zz_shift_i_6_14 = shift_i_map_36;
      6'b100101 : _zz_shift_i_6_14 = shift_i_map_37;
      6'b100110 : _zz_shift_i_6_14 = shift_i_map_38;
      6'b100111 : _zz_shift_i_6_14 = shift_i_map_39;
      6'b101000 : _zz_shift_i_6_14 = shift_i_map_40;
      6'b101001 : _zz_shift_i_6_14 = shift_i_map_41;
      6'b101010 : _zz_shift_i_6_14 = shift_i_map_42;
      6'b101011 : _zz_shift_i_6_14 = shift_i_map_43;
      6'b101100 : _zz_shift_i_6_14 = shift_i_map_44;
      6'b101101 : _zz_shift_i_6_14 = shift_i_map_45;
      6'b101110 : _zz_shift_i_6_14 = shift_i_map_46;
      6'b101111 : _zz_shift_i_6_14 = shift_i_map_47;
      6'b110000 : _zz_shift_i_6_14 = shift_i_map_48;
      6'b110001 : _zz_shift_i_6_14 = shift_i_map_49;
      6'b110010 : _zz_shift_i_6_14 = shift_i_map_50;
      6'b110011 : _zz_shift_i_6_14 = shift_i_map_51;
      6'b110100 : _zz_shift_i_6_14 = shift_i_map_52;
      6'b110101 : _zz_shift_i_6_14 = shift_i_map_53;
      6'b110110 : _zz_shift_i_6_14 = shift_i_map_54;
      6'b110111 : _zz_shift_i_6_14 = shift_i_map_55;
      6'b111000 : _zz_shift_i_6_14 = shift_i_map_56;
      6'b111001 : _zz_shift_i_6_14 = shift_i_map_57;
      6'b111010 : _zz_shift_i_6_14 = shift_i_map_58;
      6'b111011 : _zz_shift_i_6_14 = shift_i_map_59;
      6'b111100 : _zz_shift_i_6_14 = shift_i_map_60;
      6'b111101 : _zz_shift_i_6_14 = shift_i_map_61;
      6'b111110 : _zz_shift_i_6_14 = shift_i_map_62;
      default : _zz_shift_i_6_14 = shift_i_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_6_15)
      6'b000000 : _zz_shift_q_6_14 = shift_q_map_0;
      6'b000001 : _zz_shift_q_6_14 = shift_q_map_1;
      6'b000010 : _zz_shift_q_6_14 = shift_q_map_2;
      6'b000011 : _zz_shift_q_6_14 = shift_q_map_3;
      6'b000100 : _zz_shift_q_6_14 = shift_q_map_4;
      6'b000101 : _zz_shift_q_6_14 = shift_q_map_5;
      6'b000110 : _zz_shift_q_6_14 = shift_q_map_6;
      6'b000111 : _zz_shift_q_6_14 = shift_q_map_7;
      6'b001000 : _zz_shift_q_6_14 = shift_q_map_8;
      6'b001001 : _zz_shift_q_6_14 = shift_q_map_9;
      6'b001010 : _zz_shift_q_6_14 = shift_q_map_10;
      6'b001011 : _zz_shift_q_6_14 = shift_q_map_11;
      6'b001100 : _zz_shift_q_6_14 = shift_q_map_12;
      6'b001101 : _zz_shift_q_6_14 = shift_q_map_13;
      6'b001110 : _zz_shift_q_6_14 = shift_q_map_14;
      6'b001111 : _zz_shift_q_6_14 = shift_q_map_15;
      6'b010000 : _zz_shift_q_6_14 = shift_q_map_16;
      6'b010001 : _zz_shift_q_6_14 = shift_q_map_17;
      6'b010010 : _zz_shift_q_6_14 = shift_q_map_18;
      6'b010011 : _zz_shift_q_6_14 = shift_q_map_19;
      6'b010100 : _zz_shift_q_6_14 = shift_q_map_20;
      6'b010101 : _zz_shift_q_6_14 = shift_q_map_21;
      6'b010110 : _zz_shift_q_6_14 = shift_q_map_22;
      6'b010111 : _zz_shift_q_6_14 = shift_q_map_23;
      6'b011000 : _zz_shift_q_6_14 = shift_q_map_24;
      6'b011001 : _zz_shift_q_6_14 = shift_q_map_25;
      6'b011010 : _zz_shift_q_6_14 = shift_q_map_26;
      6'b011011 : _zz_shift_q_6_14 = shift_q_map_27;
      6'b011100 : _zz_shift_q_6_14 = shift_q_map_28;
      6'b011101 : _zz_shift_q_6_14 = shift_q_map_29;
      6'b011110 : _zz_shift_q_6_14 = shift_q_map_30;
      6'b011111 : _zz_shift_q_6_14 = shift_q_map_31;
      6'b100000 : _zz_shift_q_6_14 = shift_q_map_32;
      6'b100001 : _zz_shift_q_6_14 = shift_q_map_33;
      6'b100010 : _zz_shift_q_6_14 = shift_q_map_34;
      6'b100011 : _zz_shift_q_6_14 = shift_q_map_35;
      6'b100100 : _zz_shift_q_6_14 = shift_q_map_36;
      6'b100101 : _zz_shift_q_6_14 = shift_q_map_37;
      6'b100110 : _zz_shift_q_6_14 = shift_q_map_38;
      6'b100111 : _zz_shift_q_6_14 = shift_q_map_39;
      6'b101000 : _zz_shift_q_6_14 = shift_q_map_40;
      6'b101001 : _zz_shift_q_6_14 = shift_q_map_41;
      6'b101010 : _zz_shift_q_6_14 = shift_q_map_42;
      6'b101011 : _zz_shift_q_6_14 = shift_q_map_43;
      6'b101100 : _zz_shift_q_6_14 = shift_q_map_44;
      6'b101101 : _zz_shift_q_6_14 = shift_q_map_45;
      6'b101110 : _zz_shift_q_6_14 = shift_q_map_46;
      6'b101111 : _zz_shift_q_6_14 = shift_q_map_47;
      6'b110000 : _zz_shift_q_6_14 = shift_q_map_48;
      6'b110001 : _zz_shift_q_6_14 = shift_q_map_49;
      6'b110010 : _zz_shift_q_6_14 = shift_q_map_50;
      6'b110011 : _zz_shift_q_6_14 = shift_q_map_51;
      6'b110100 : _zz_shift_q_6_14 = shift_q_map_52;
      6'b110101 : _zz_shift_q_6_14 = shift_q_map_53;
      6'b110110 : _zz_shift_q_6_14 = shift_q_map_54;
      6'b110111 : _zz_shift_q_6_14 = shift_q_map_55;
      6'b111000 : _zz_shift_q_6_14 = shift_q_map_56;
      6'b111001 : _zz_shift_q_6_14 = shift_q_map_57;
      6'b111010 : _zz_shift_q_6_14 = shift_q_map_58;
      6'b111011 : _zz_shift_q_6_14 = shift_q_map_59;
      6'b111100 : _zz_shift_q_6_14 = shift_q_map_60;
      6'b111101 : _zz_shift_q_6_14 = shift_q_map_61;
      6'b111110 : _zz_shift_q_6_14 = shift_q_map_62;
      default : _zz_shift_q_6_14 = shift_q_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_7_15)
      6'b000000 : _zz_shift_i_7_14 = shift_i_map_0;
      6'b000001 : _zz_shift_i_7_14 = shift_i_map_1;
      6'b000010 : _zz_shift_i_7_14 = shift_i_map_2;
      6'b000011 : _zz_shift_i_7_14 = shift_i_map_3;
      6'b000100 : _zz_shift_i_7_14 = shift_i_map_4;
      6'b000101 : _zz_shift_i_7_14 = shift_i_map_5;
      6'b000110 : _zz_shift_i_7_14 = shift_i_map_6;
      6'b000111 : _zz_shift_i_7_14 = shift_i_map_7;
      6'b001000 : _zz_shift_i_7_14 = shift_i_map_8;
      6'b001001 : _zz_shift_i_7_14 = shift_i_map_9;
      6'b001010 : _zz_shift_i_7_14 = shift_i_map_10;
      6'b001011 : _zz_shift_i_7_14 = shift_i_map_11;
      6'b001100 : _zz_shift_i_7_14 = shift_i_map_12;
      6'b001101 : _zz_shift_i_7_14 = shift_i_map_13;
      6'b001110 : _zz_shift_i_7_14 = shift_i_map_14;
      6'b001111 : _zz_shift_i_7_14 = shift_i_map_15;
      6'b010000 : _zz_shift_i_7_14 = shift_i_map_16;
      6'b010001 : _zz_shift_i_7_14 = shift_i_map_17;
      6'b010010 : _zz_shift_i_7_14 = shift_i_map_18;
      6'b010011 : _zz_shift_i_7_14 = shift_i_map_19;
      6'b010100 : _zz_shift_i_7_14 = shift_i_map_20;
      6'b010101 : _zz_shift_i_7_14 = shift_i_map_21;
      6'b010110 : _zz_shift_i_7_14 = shift_i_map_22;
      6'b010111 : _zz_shift_i_7_14 = shift_i_map_23;
      6'b011000 : _zz_shift_i_7_14 = shift_i_map_24;
      6'b011001 : _zz_shift_i_7_14 = shift_i_map_25;
      6'b011010 : _zz_shift_i_7_14 = shift_i_map_26;
      6'b011011 : _zz_shift_i_7_14 = shift_i_map_27;
      6'b011100 : _zz_shift_i_7_14 = shift_i_map_28;
      6'b011101 : _zz_shift_i_7_14 = shift_i_map_29;
      6'b011110 : _zz_shift_i_7_14 = shift_i_map_30;
      6'b011111 : _zz_shift_i_7_14 = shift_i_map_31;
      6'b100000 : _zz_shift_i_7_14 = shift_i_map_32;
      6'b100001 : _zz_shift_i_7_14 = shift_i_map_33;
      6'b100010 : _zz_shift_i_7_14 = shift_i_map_34;
      6'b100011 : _zz_shift_i_7_14 = shift_i_map_35;
      6'b100100 : _zz_shift_i_7_14 = shift_i_map_36;
      6'b100101 : _zz_shift_i_7_14 = shift_i_map_37;
      6'b100110 : _zz_shift_i_7_14 = shift_i_map_38;
      6'b100111 : _zz_shift_i_7_14 = shift_i_map_39;
      6'b101000 : _zz_shift_i_7_14 = shift_i_map_40;
      6'b101001 : _zz_shift_i_7_14 = shift_i_map_41;
      6'b101010 : _zz_shift_i_7_14 = shift_i_map_42;
      6'b101011 : _zz_shift_i_7_14 = shift_i_map_43;
      6'b101100 : _zz_shift_i_7_14 = shift_i_map_44;
      6'b101101 : _zz_shift_i_7_14 = shift_i_map_45;
      6'b101110 : _zz_shift_i_7_14 = shift_i_map_46;
      6'b101111 : _zz_shift_i_7_14 = shift_i_map_47;
      6'b110000 : _zz_shift_i_7_14 = shift_i_map_48;
      6'b110001 : _zz_shift_i_7_14 = shift_i_map_49;
      6'b110010 : _zz_shift_i_7_14 = shift_i_map_50;
      6'b110011 : _zz_shift_i_7_14 = shift_i_map_51;
      6'b110100 : _zz_shift_i_7_14 = shift_i_map_52;
      6'b110101 : _zz_shift_i_7_14 = shift_i_map_53;
      6'b110110 : _zz_shift_i_7_14 = shift_i_map_54;
      6'b110111 : _zz_shift_i_7_14 = shift_i_map_55;
      6'b111000 : _zz_shift_i_7_14 = shift_i_map_56;
      6'b111001 : _zz_shift_i_7_14 = shift_i_map_57;
      6'b111010 : _zz_shift_i_7_14 = shift_i_map_58;
      6'b111011 : _zz_shift_i_7_14 = shift_i_map_59;
      6'b111100 : _zz_shift_i_7_14 = shift_i_map_60;
      6'b111101 : _zz_shift_i_7_14 = shift_i_map_61;
      6'b111110 : _zz_shift_i_7_14 = shift_i_map_62;
      default : _zz_shift_i_7_14 = shift_i_map_63;
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_7_15)
      6'b000000 : _zz_shift_q_7_14 = shift_q_map_0;
      6'b000001 : _zz_shift_q_7_14 = shift_q_map_1;
      6'b000010 : _zz_shift_q_7_14 = shift_q_map_2;
      6'b000011 : _zz_shift_q_7_14 = shift_q_map_3;
      6'b000100 : _zz_shift_q_7_14 = shift_q_map_4;
      6'b000101 : _zz_shift_q_7_14 = shift_q_map_5;
      6'b000110 : _zz_shift_q_7_14 = shift_q_map_6;
      6'b000111 : _zz_shift_q_7_14 = shift_q_map_7;
      6'b001000 : _zz_shift_q_7_14 = shift_q_map_8;
      6'b001001 : _zz_shift_q_7_14 = shift_q_map_9;
      6'b001010 : _zz_shift_q_7_14 = shift_q_map_10;
      6'b001011 : _zz_shift_q_7_14 = shift_q_map_11;
      6'b001100 : _zz_shift_q_7_14 = shift_q_map_12;
      6'b001101 : _zz_shift_q_7_14 = shift_q_map_13;
      6'b001110 : _zz_shift_q_7_14 = shift_q_map_14;
      6'b001111 : _zz_shift_q_7_14 = shift_q_map_15;
      6'b010000 : _zz_shift_q_7_14 = shift_q_map_16;
      6'b010001 : _zz_shift_q_7_14 = shift_q_map_17;
      6'b010010 : _zz_shift_q_7_14 = shift_q_map_18;
      6'b010011 : _zz_shift_q_7_14 = shift_q_map_19;
      6'b010100 : _zz_shift_q_7_14 = shift_q_map_20;
      6'b010101 : _zz_shift_q_7_14 = shift_q_map_21;
      6'b010110 : _zz_shift_q_7_14 = shift_q_map_22;
      6'b010111 : _zz_shift_q_7_14 = shift_q_map_23;
      6'b011000 : _zz_shift_q_7_14 = shift_q_map_24;
      6'b011001 : _zz_shift_q_7_14 = shift_q_map_25;
      6'b011010 : _zz_shift_q_7_14 = shift_q_map_26;
      6'b011011 : _zz_shift_q_7_14 = shift_q_map_27;
      6'b011100 : _zz_shift_q_7_14 = shift_q_map_28;
      6'b011101 : _zz_shift_q_7_14 = shift_q_map_29;
      6'b011110 : _zz_shift_q_7_14 = shift_q_map_30;
      6'b011111 : _zz_shift_q_7_14 = shift_q_map_31;
      6'b100000 : _zz_shift_q_7_14 = shift_q_map_32;
      6'b100001 : _zz_shift_q_7_14 = shift_q_map_33;
      6'b100010 : _zz_shift_q_7_14 = shift_q_map_34;
      6'b100011 : _zz_shift_q_7_14 = shift_q_map_35;
      6'b100100 : _zz_shift_q_7_14 = shift_q_map_36;
      6'b100101 : _zz_shift_q_7_14 = shift_q_map_37;
      6'b100110 : _zz_shift_q_7_14 = shift_q_map_38;
      6'b100111 : _zz_shift_q_7_14 = shift_q_map_39;
      6'b101000 : _zz_shift_q_7_14 = shift_q_map_40;
      6'b101001 : _zz_shift_q_7_14 = shift_q_map_41;
      6'b101010 : _zz_shift_q_7_14 = shift_q_map_42;
      6'b101011 : _zz_shift_q_7_14 = shift_q_map_43;
      6'b101100 : _zz_shift_q_7_14 = shift_q_map_44;
      6'b101101 : _zz_shift_q_7_14 = shift_q_map_45;
      6'b101110 : _zz_shift_q_7_14 = shift_q_map_46;
      6'b101111 : _zz_shift_q_7_14 = shift_q_map_47;
      6'b110000 : _zz_shift_q_7_14 = shift_q_map_48;
      6'b110001 : _zz_shift_q_7_14 = shift_q_map_49;
      6'b110010 : _zz_shift_q_7_14 = shift_q_map_50;
      6'b110011 : _zz_shift_q_7_14 = shift_q_map_51;
      6'b110100 : _zz_shift_q_7_14 = shift_q_map_52;
      6'b110101 : _zz_shift_q_7_14 = shift_q_map_53;
      6'b110110 : _zz_shift_q_7_14 = shift_q_map_54;
      6'b110111 : _zz_shift_q_7_14 = shift_q_map_55;
      6'b111000 : _zz_shift_q_7_14 = shift_q_map_56;
      6'b111001 : _zz_shift_q_7_14 = shift_q_map_57;
      6'b111010 : _zz_shift_q_7_14 = shift_q_map_58;
      6'b111011 : _zz_shift_q_7_14 = shift_q_map_59;
      6'b111100 : _zz_shift_q_7_14 = shift_q_map_60;
      6'b111101 : _zz_shift_q_7_14 = shift_q_map_61;
      6'b111110 : _zz_shift_q_7_14 = shift_q_map_62;
      default : _zz_shift_q_7_14 = shift_q_map_63;
    endcase
  end

  assign _zz_1 = ({63'd0,1'b1} <<< w_addr);
  assign _zz_2 = ({63'd0,1'b1} <<< w_addr);
  assign base_sub_iqs_payload_0_cha_i = mIMOReceiverUnit_8_base_sub_iq_payload_cha_i;
  assign base_sub_iqs_payload_0_cha_q = mIMOReceiverUnit_8_base_sub_iq_payload_cha_q;
  assign base_sub_valid_vec_0 = mIMOReceiverUnit_8_base_sub_iq_valid;
  assign mIMOReceiverUnit_8_shift_i_0 = _zz_shift_i_0;
  assign mIMOReceiverUnit_8_shift_q_0 = _zz_shift_q_0;
  assign mIMOReceiverUnit_8_shift_i_1 = _zz_shift_i_1;
  assign mIMOReceiverUnit_8_shift_q_1 = _zz_shift_q_1;
  assign mIMOReceiverUnit_8_shift_i_2 = _zz_shift_i_2;
  assign mIMOReceiverUnit_8_shift_q_2 = _zz_shift_q_2;
  assign mIMOReceiverUnit_8_shift_i_3 = _zz_shift_i_3;
  assign mIMOReceiverUnit_8_shift_q_3 = _zz_shift_q_3;
  assign mIMOReceiverUnit_8_shift_i_4 = _zz_shift_i_4;
  assign mIMOReceiverUnit_8_shift_q_4 = _zz_shift_q_4;
  assign mIMOReceiverUnit_8_shift_i_5 = _zz_shift_i_5;
  assign mIMOReceiverUnit_8_shift_q_5 = _zz_shift_q_5;
  assign mIMOReceiverUnit_8_shift_i_6 = _zz_shift_i_6;
  assign mIMOReceiverUnit_8_shift_q_6 = _zz_shift_q_6;
  assign mIMOReceiverUnit_8_shift_i_7 = _zz_shift_i_7;
  assign mIMOReceiverUnit_8_shift_q_7 = _zz_shift_q_7;
  assign base_sub_iqs_payload_1_cha_i = mIMOReceiverUnit_9_base_sub_iq_payload_cha_i;
  assign base_sub_iqs_payload_1_cha_q = mIMOReceiverUnit_9_base_sub_iq_payload_cha_q;
  assign base_sub_valid_vec_1 = mIMOReceiverUnit_9_base_sub_iq_valid;
  assign mIMOReceiverUnit_9_shift_i_0 = _zz_shift_i_0_2;
  assign mIMOReceiverUnit_9_shift_q_0 = _zz_shift_q_0_2;
  assign mIMOReceiverUnit_9_shift_i_1 = _zz_shift_i_1_2;
  assign mIMOReceiverUnit_9_shift_q_1 = _zz_shift_q_1_2;
  assign mIMOReceiverUnit_9_shift_i_2 = _zz_shift_i_2_2;
  assign mIMOReceiverUnit_9_shift_q_2 = _zz_shift_q_2_2;
  assign mIMOReceiverUnit_9_shift_i_3 = _zz_shift_i_3_2;
  assign mIMOReceiverUnit_9_shift_q_3 = _zz_shift_q_3_2;
  assign mIMOReceiverUnit_9_shift_i_4 = _zz_shift_i_4_2;
  assign mIMOReceiverUnit_9_shift_q_4 = _zz_shift_q_4_2;
  assign mIMOReceiverUnit_9_shift_i_5 = _zz_shift_i_5_2;
  assign mIMOReceiverUnit_9_shift_q_5 = _zz_shift_q_5_2;
  assign mIMOReceiverUnit_9_shift_i_6 = _zz_shift_i_6_2;
  assign mIMOReceiverUnit_9_shift_q_6 = _zz_shift_q_6_2;
  assign mIMOReceiverUnit_9_shift_i_7 = _zz_shift_i_7_2;
  assign mIMOReceiverUnit_9_shift_q_7 = _zz_shift_q_7_2;
  assign base_sub_iqs_payload_2_cha_i = mIMOReceiverUnit_10_base_sub_iq_payload_cha_i;
  assign base_sub_iqs_payload_2_cha_q = mIMOReceiverUnit_10_base_sub_iq_payload_cha_q;
  assign base_sub_valid_vec_2 = mIMOReceiverUnit_10_base_sub_iq_valid;
  assign mIMOReceiverUnit_10_shift_i_0 = _zz_shift_i_0_4;
  assign mIMOReceiverUnit_10_shift_q_0 = _zz_shift_q_0_4;
  assign mIMOReceiverUnit_10_shift_i_1 = _zz_shift_i_1_4;
  assign mIMOReceiverUnit_10_shift_q_1 = _zz_shift_q_1_4;
  assign mIMOReceiverUnit_10_shift_i_2 = _zz_shift_i_2_4;
  assign mIMOReceiverUnit_10_shift_q_2 = _zz_shift_q_2_4;
  assign mIMOReceiverUnit_10_shift_i_3 = _zz_shift_i_3_4;
  assign mIMOReceiverUnit_10_shift_q_3 = _zz_shift_q_3_4;
  assign mIMOReceiverUnit_10_shift_i_4 = _zz_shift_i_4_4;
  assign mIMOReceiverUnit_10_shift_q_4 = _zz_shift_q_4_4;
  assign mIMOReceiverUnit_10_shift_i_5 = _zz_shift_i_5_4;
  assign mIMOReceiverUnit_10_shift_q_5 = _zz_shift_q_5_4;
  assign mIMOReceiverUnit_10_shift_i_6 = _zz_shift_i_6_4;
  assign mIMOReceiverUnit_10_shift_q_6 = _zz_shift_q_6_4;
  assign mIMOReceiverUnit_10_shift_i_7 = _zz_shift_i_7_4;
  assign mIMOReceiverUnit_10_shift_q_7 = _zz_shift_q_7_4;
  assign base_sub_iqs_payload_3_cha_i = mIMOReceiverUnit_11_base_sub_iq_payload_cha_i;
  assign base_sub_iqs_payload_3_cha_q = mIMOReceiverUnit_11_base_sub_iq_payload_cha_q;
  assign base_sub_valid_vec_3 = mIMOReceiverUnit_11_base_sub_iq_valid;
  assign mIMOReceiverUnit_11_shift_i_0 = _zz_shift_i_0_6;
  assign mIMOReceiverUnit_11_shift_q_0 = _zz_shift_q_0_6;
  assign mIMOReceiverUnit_11_shift_i_1 = _zz_shift_i_1_6;
  assign mIMOReceiverUnit_11_shift_q_1 = _zz_shift_q_1_6;
  assign mIMOReceiverUnit_11_shift_i_2 = _zz_shift_i_2_6;
  assign mIMOReceiverUnit_11_shift_q_2 = _zz_shift_q_2_6;
  assign mIMOReceiverUnit_11_shift_i_3 = _zz_shift_i_3_6;
  assign mIMOReceiverUnit_11_shift_q_3 = _zz_shift_q_3_6;
  assign mIMOReceiverUnit_11_shift_i_4 = _zz_shift_i_4_6;
  assign mIMOReceiverUnit_11_shift_q_4 = _zz_shift_q_4_6;
  assign mIMOReceiverUnit_11_shift_i_5 = _zz_shift_i_5_6;
  assign mIMOReceiverUnit_11_shift_q_5 = _zz_shift_q_5_6;
  assign mIMOReceiverUnit_11_shift_i_6 = _zz_shift_i_6_6;
  assign mIMOReceiverUnit_11_shift_q_6 = _zz_shift_q_6_6;
  assign mIMOReceiverUnit_11_shift_i_7 = _zz_shift_i_7_6;
  assign mIMOReceiverUnit_11_shift_q_7 = _zz_shift_q_7_6;
  assign base_sub_iqs_payload_4_cha_i = mIMOReceiverUnit_12_base_sub_iq_payload_cha_i;
  assign base_sub_iqs_payload_4_cha_q = mIMOReceiverUnit_12_base_sub_iq_payload_cha_q;
  assign base_sub_valid_vec_4 = mIMOReceiverUnit_12_base_sub_iq_valid;
  assign mIMOReceiverUnit_12_shift_i_0 = _zz_shift_i_0_8;
  assign mIMOReceiverUnit_12_shift_q_0 = _zz_shift_q_0_8;
  assign mIMOReceiverUnit_12_shift_i_1 = _zz_shift_i_1_8;
  assign mIMOReceiverUnit_12_shift_q_1 = _zz_shift_q_1_8;
  assign mIMOReceiverUnit_12_shift_i_2 = _zz_shift_i_2_8;
  assign mIMOReceiverUnit_12_shift_q_2 = _zz_shift_q_2_8;
  assign mIMOReceiverUnit_12_shift_i_3 = _zz_shift_i_3_8;
  assign mIMOReceiverUnit_12_shift_q_3 = _zz_shift_q_3_8;
  assign mIMOReceiverUnit_12_shift_i_4 = _zz_shift_i_4_8;
  assign mIMOReceiverUnit_12_shift_q_4 = _zz_shift_q_4_8;
  assign mIMOReceiverUnit_12_shift_i_5 = _zz_shift_i_5_8;
  assign mIMOReceiverUnit_12_shift_q_5 = _zz_shift_q_5_8;
  assign mIMOReceiverUnit_12_shift_i_6 = _zz_shift_i_6_8;
  assign mIMOReceiverUnit_12_shift_q_6 = _zz_shift_q_6_8;
  assign mIMOReceiverUnit_12_shift_i_7 = _zz_shift_i_7_8;
  assign mIMOReceiverUnit_12_shift_q_7 = _zz_shift_q_7_8;
  assign base_sub_iqs_payload_5_cha_i = mIMOReceiverUnit_13_base_sub_iq_payload_cha_i;
  assign base_sub_iqs_payload_5_cha_q = mIMOReceiverUnit_13_base_sub_iq_payload_cha_q;
  assign base_sub_valid_vec_5 = mIMOReceiverUnit_13_base_sub_iq_valid;
  assign mIMOReceiverUnit_13_shift_i_0 = _zz_shift_i_0_10;
  assign mIMOReceiverUnit_13_shift_q_0 = _zz_shift_q_0_10;
  assign mIMOReceiverUnit_13_shift_i_1 = _zz_shift_i_1_10;
  assign mIMOReceiverUnit_13_shift_q_1 = _zz_shift_q_1_10;
  assign mIMOReceiverUnit_13_shift_i_2 = _zz_shift_i_2_10;
  assign mIMOReceiverUnit_13_shift_q_2 = _zz_shift_q_2_10;
  assign mIMOReceiverUnit_13_shift_i_3 = _zz_shift_i_3_10;
  assign mIMOReceiverUnit_13_shift_q_3 = _zz_shift_q_3_10;
  assign mIMOReceiverUnit_13_shift_i_4 = _zz_shift_i_4_10;
  assign mIMOReceiverUnit_13_shift_q_4 = _zz_shift_q_4_10;
  assign mIMOReceiverUnit_13_shift_i_5 = _zz_shift_i_5_10;
  assign mIMOReceiverUnit_13_shift_q_5 = _zz_shift_q_5_10;
  assign mIMOReceiverUnit_13_shift_i_6 = _zz_shift_i_6_10;
  assign mIMOReceiverUnit_13_shift_q_6 = _zz_shift_q_6_10;
  assign mIMOReceiverUnit_13_shift_i_7 = _zz_shift_i_7_10;
  assign mIMOReceiverUnit_13_shift_q_7 = _zz_shift_q_7_10;
  assign base_sub_iqs_payload_6_cha_i = mIMOReceiverUnit_14_base_sub_iq_payload_cha_i;
  assign base_sub_iqs_payload_6_cha_q = mIMOReceiverUnit_14_base_sub_iq_payload_cha_q;
  assign base_sub_valid_vec_6 = mIMOReceiverUnit_14_base_sub_iq_valid;
  assign mIMOReceiverUnit_14_shift_i_0 = _zz_shift_i_0_12;
  assign mIMOReceiverUnit_14_shift_q_0 = _zz_shift_q_0_12;
  assign mIMOReceiverUnit_14_shift_i_1 = _zz_shift_i_1_12;
  assign mIMOReceiverUnit_14_shift_q_1 = _zz_shift_q_1_12;
  assign mIMOReceiverUnit_14_shift_i_2 = _zz_shift_i_2_12;
  assign mIMOReceiverUnit_14_shift_q_2 = _zz_shift_q_2_12;
  assign mIMOReceiverUnit_14_shift_i_3 = _zz_shift_i_3_12;
  assign mIMOReceiverUnit_14_shift_q_3 = _zz_shift_q_3_12;
  assign mIMOReceiverUnit_14_shift_i_4 = _zz_shift_i_4_12;
  assign mIMOReceiverUnit_14_shift_q_4 = _zz_shift_q_4_12;
  assign mIMOReceiverUnit_14_shift_i_5 = _zz_shift_i_5_12;
  assign mIMOReceiverUnit_14_shift_q_5 = _zz_shift_q_5_12;
  assign mIMOReceiverUnit_14_shift_i_6 = _zz_shift_i_6_12;
  assign mIMOReceiverUnit_14_shift_q_6 = _zz_shift_q_6_12;
  assign mIMOReceiverUnit_14_shift_i_7 = _zz_shift_i_7_12;
  assign mIMOReceiverUnit_14_shift_q_7 = _zz_shift_q_7_12;
  assign base_sub_iqs_payload_7_cha_i = mIMOReceiverUnit_15_base_sub_iq_payload_cha_i;
  assign base_sub_iqs_payload_7_cha_q = mIMOReceiverUnit_15_base_sub_iq_payload_cha_q;
  assign base_sub_valid_vec_7 = mIMOReceiverUnit_15_base_sub_iq_valid;
  assign mIMOReceiverUnit_15_shift_i_0 = _zz_shift_i_0_14;
  assign mIMOReceiverUnit_15_shift_q_0 = _zz_shift_q_0_14;
  assign mIMOReceiverUnit_15_shift_i_1 = _zz_shift_i_1_14;
  assign mIMOReceiverUnit_15_shift_q_1 = _zz_shift_q_1_14;
  assign mIMOReceiverUnit_15_shift_i_2 = _zz_shift_i_2_14;
  assign mIMOReceiverUnit_15_shift_q_2 = _zz_shift_q_2_14;
  assign mIMOReceiverUnit_15_shift_i_3 = _zz_shift_i_3_14;
  assign mIMOReceiverUnit_15_shift_q_3 = _zz_shift_q_3_14;
  assign mIMOReceiverUnit_15_shift_i_4 = _zz_shift_i_4_14;
  assign mIMOReceiverUnit_15_shift_q_4 = _zz_shift_q_4_14;
  assign mIMOReceiverUnit_15_shift_i_5 = _zz_shift_i_5_14;
  assign mIMOReceiverUnit_15_shift_q_5 = _zz_shift_q_5_14;
  assign mIMOReceiverUnit_15_shift_i_6 = _zz_shift_i_6_14;
  assign mIMOReceiverUnit_15_shift_q_6 = _zz_shift_q_6_14;
  assign mIMOReceiverUnit_15_shift_i_7 = _zz_shift_i_7_14;
  assign mIMOReceiverUnit_15_shift_q_7 = _zz_shift_q_7_14;
  assign base_sub_iqs_valid = (((((((base_sub_valid_vec_0 && base_sub_valid_vec_1) && base_sub_valid_vec_2) && base_sub_valid_vec_3) && base_sub_valid_vec_4) && base_sub_valid_vec_5) && base_sub_valid_vec_6) && base_sub_valid_vec_7);
  assign mod_iq_ready = (! w_en);
  always @(posedge rf_clk) begin
    if(w_en) begin
      if(w_sel) begin
        if(_zz_1[0]) begin
          shift_i_map_0 <= w_data;
        end
        if(_zz_1[1]) begin
          shift_i_map_1 <= w_data;
        end
        if(_zz_1[2]) begin
          shift_i_map_2 <= w_data;
        end
        if(_zz_1[3]) begin
          shift_i_map_3 <= w_data;
        end
        if(_zz_1[4]) begin
          shift_i_map_4 <= w_data;
        end
        if(_zz_1[5]) begin
          shift_i_map_5 <= w_data;
        end
        if(_zz_1[6]) begin
          shift_i_map_6 <= w_data;
        end
        if(_zz_1[7]) begin
          shift_i_map_7 <= w_data;
        end
        if(_zz_1[8]) begin
          shift_i_map_8 <= w_data;
        end
        if(_zz_1[9]) begin
          shift_i_map_9 <= w_data;
        end
        if(_zz_1[10]) begin
          shift_i_map_10 <= w_data;
        end
        if(_zz_1[11]) begin
          shift_i_map_11 <= w_data;
        end
        if(_zz_1[12]) begin
          shift_i_map_12 <= w_data;
        end
        if(_zz_1[13]) begin
          shift_i_map_13 <= w_data;
        end
        if(_zz_1[14]) begin
          shift_i_map_14 <= w_data;
        end
        if(_zz_1[15]) begin
          shift_i_map_15 <= w_data;
        end
        if(_zz_1[16]) begin
          shift_i_map_16 <= w_data;
        end
        if(_zz_1[17]) begin
          shift_i_map_17 <= w_data;
        end
        if(_zz_1[18]) begin
          shift_i_map_18 <= w_data;
        end
        if(_zz_1[19]) begin
          shift_i_map_19 <= w_data;
        end
        if(_zz_1[20]) begin
          shift_i_map_20 <= w_data;
        end
        if(_zz_1[21]) begin
          shift_i_map_21 <= w_data;
        end
        if(_zz_1[22]) begin
          shift_i_map_22 <= w_data;
        end
        if(_zz_1[23]) begin
          shift_i_map_23 <= w_data;
        end
        if(_zz_1[24]) begin
          shift_i_map_24 <= w_data;
        end
        if(_zz_1[25]) begin
          shift_i_map_25 <= w_data;
        end
        if(_zz_1[26]) begin
          shift_i_map_26 <= w_data;
        end
        if(_zz_1[27]) begin
          shift_i_map_27 <= w_data;
        end
        if(_zz_1[28]) begin
          shift_i_map_28 <= w_data;
        end
        if(_zz_1[29]) begin
          shift_i_map_29 <= w_data;
        end
        if(_zz_1[30]) begin
          shift_i_map_30 <= w_data;
        end
        if(_zz_1[31]) begin
          shift_i_map_31 <= w_data;
        end
        if(_zz_1[32]) begin
          shift_i_map_32 <= w_data;
        end
        if(_zz_1[33]) begin
          shift_i_map_33 <= w_data;
        end
        if(_zz_1[34]) begin
          shift_i_map_34 <= w_data;
        end
        if(_zz_1[35]) begin
          shift_i_map_35 <= w_data;
        end
        if(_zz_1[36]) begin
          shift_i_map_36 <= w_data;
        end
        if(_zz_1[37]) begin
          shift_i_map_37 <= w_data;
        end
        if(_zz_1[38]) begin
          shift_i_map_38 <= w_data;
        end
        if(_zz_1[39]) begin
          shift_i_map_39 <= w_data;
        end
        if(_zz_1[40]) begin
          shift_i_map_40 <= w_data;
        end
        if(_zz_1[41]) begin
          shift_i_map_41 <= w_data;
        end
        if(_zz_1[42]) begin
          shift_i_map_42 <= w_data;
        end
        if(_zz_1[43]) begin
          shift_i_map_43 <= w_data;
        end
        if(_zz_1[44]) begin
          shift_i_map_44 <= w_data;
        end
        if(_zz_1[45]) begin
          shift_i_map_45 <= w_data;
        end
        if(_zz_1[46]) begin
          shift_i_map_46 <= w_data;
        end
        if(_zz_1[47]) begin
          shift_i_map_47 <= w_data;
        end
        if(_zz_1[48]) begin
          shift_i_map_48 <= w_data;
        end
        if(_zz_1[49]) begin
          shift_i_map_49 <= w_data;
        end
        if(_zz_1[50]) begin
          shift_i_map_50 <= w_data;
        end
        if(_zz_1[51]) begin
          shift_i_map_51 <= w_data;
        end
        if(_zz_1[52]) begin
          shift_i_map_52 <= w_data;
        end
        if(_zz_1[53]) begin
          shift_i_map_53 <= w_data;
        end
        if(_zz_1[54]) begin
          shift_i_map_54 <= w_data;
        end
        if(_zz_1[55]) begin
          shift_i_map_55 <= w_data;
        end
        if(_zz_1[56]) begin
          shift_i_map_56 <= w_data;
        end
        if(_zz_1[57]) begin
          shift_i_map_57 <= w_data;
        end
        if(_zz_1[58]) begin
          shift_i_map_58 <= w_data;
        end
        if(_zz_1[59]) begin
          shift_i_map_59 <= w_data;
        end
        if(_zz_1[60]) begin
          shift_i_map_60 <= w_data;
        end
        if(_zz_1[61]) begin
          shift_i_map_61 <= w_data;
        end
        if(_zz_1[62]) begin
          shift_i_map_62 <= w_data;
        end
        if(_zz_1[63]) begin
          shift_i_map_63 <= w_data;
        end
      end else begin
        if(_zz_2[0]) begin
          shift_q_map_0 <= w_data;
        end
        if(_zz_2[1]) begin
          shift_q_map_1 <= w_data;
        end
        if(_zz_2[2]) begin
          shift_q_map_2 <= w_data;
        end
        if(_zz_2[3]) begin
          shift_q_map_3 <= w_data;
        end
        if(_zz_2[4]) begin
          shift_q_map_4 <= w_data;
        end
        if(_zz_2[5]) begin
          shift_q_map_5 <= w_data;
        end
        if(_zz_2[6]) begin
          shift_q_map_6 <= w_data;
        end
        if(_zz_2[7]) begin
          shift_q_map_7 <= w_data;
        end
        if(_zz_2[8]) begin
          shift_q_map_8 <= w_data;
        end
        if(_zz_2[9]) begin
          shift_q_map_9 <= w_data;
        end
        if(_zz_2[10]) begin
          shift_q_map_10 <= w_data;
        end
        if(_zz_2[11]) begin
          shift_q_map_11 <= w_data;
        end
        if(_zz_2[12]) begin
          shift_q_map_12 <= w_data;
        end
        if(_zz_2[13]) begin
          shift_q_map_13 <= w_data;
        end
        if(_zz_2[14]) begin
          shift_q_map_14 <= w_data;
        end
        if(_zz_2[15]) begin
          shift_q_map_15 <= w_data;
        end
        if(_zz_2[16]) begin
          shift_q_map_16 <= w_data;
        end
        if(_zz_2[17]) begin
          shift_q_map_17 <= w_data;
        end
        if(_zz_2[18]) begin
          shift_q_map_18 <= w_data;
        end
        if(_zz_2[19]) begin
          shift_q_map_19 <= w_data;
        end
        if(_zz_2[20]) begin
          shift_q_map_20 <= w_data;
        end
        if(_zz_2[21]) begin
          shift_q_map_21 <= w_data;
        end
        if(_zz_2[22]) begin
          shift_q_map_22 <= w_data;
        end
        if(_zz_2[23]) begin
          shift_q_map_23 <= w_data;
        end
        if(_zz_2[24]) begin
          shift_q_map_24 <= w_data;
        end
        if(_zz_2[25]) begin
          shift_q_map_25 <= w_data;
        end
        if(_zz_2[26]) begin
          shift_q_map_26 <= w_data;
        end
        if(_zz_2[27]) begin
          shift_q_map_27 <= w_data;
        end
        if(_zz_2[28]) begin
          shift_q_map_28 <= w_data;
        end
        if(_zz_2[29]) begin
          shift_q_map_29 <= w_data;
        end
        if(_zz_2[30]) begin
          shift_q_map_30 <= w_data;
        end
        if(_zz_2[31]) begin
          shift_q_map_31 <= w_data;
        end
        if(_zz_2[32]) begin
          shift_q_map_32 <= w_data;
        end
        if(_zz_2[33]) begin
          shift_q_map_33 <= w_data;
        end
        if(_zz_2[34]) begin
          shift_q_map_34 <= w_data;
        end
        if(_zz_2[35]) begin
          shift_q_map_35 <= w_data;
        end
        if(_zz_2[36]) begin
          shift_q_map_36 <= w_data;
        end
        if(_zz_2[37]) begin
          shift_q_map_37 <= w_data;
        end
        if(_zz_2[38]) begin
          shift_q_map_38 <= w_data;
        end
        if(_zz_2[39]) begin
          shift_q_map_39 <= w_data;
        end
        if(_zz_2[40]) begin
          shift_q_map_40 <= w_data;
        end
        if(_zz_2[41]) begin
          shift_q_map_41 <= w_data;
        end
        if(_zz_2[42]) begin
          shift_q_map_42 <= w_data;
        end
        if(_zz_2[43]) begin
          shift_q_map_43 <= w_data;
        end
        if(_zz_2[44]) begin
          shift_q_map_44 <= w_data;
        end
        if(_zz_2[45]) begin
          shift_q_map_45 <= w_data;
        end
        if(_zz_2[46]) begin
          shift_q_map_46 <= w_data;
        end
        if(_zz_2[47]) begin
          shift_q_map_47 <= w_data;
        end
        if(_zz_2[48]) begin
          shift_q_map_48 <= w_data;
        end
        if(_zz_2[49]) begin
          shift_q_map_49 <= w_data;
        end
        if(_zz_2[50]) begin
          shift_q_map_50 <= w_data;
        end
        if(_zz_2[51]) begin
          shift_q_map_51 <= w_data;
        end
        if(_zz_2[52]) begin
          shift_q_map_52 <= w_data;
        end
        if(_zz_2[53]) begin
          shift_q_map_53 <= w_data;
        end
        if(_zz_2[54]) begin
          shift_q_map_54 <= w_data;
        end
        if(_zz_2[55]) begin
          shift_q_map_55 <= w_data;
        end
        if(_zz_2[56]) begin
          shift_q_map_56 <= w_data;
        end
        if(_zz_2[57]) begin
          shift_q_map_57 <= w_data;
        end
        if(_zz_2[58]) begin
          shift_q_map_58 <= w_data;
        end
        if(_zz_2[59]) begin
          shift_q_map_59 <= w_data;
        end
        if(_zz_2[60]) begin
          shift_q_map_60 <= w_data;
        end
        if(_zz_2[61]) begin
          shift_q_map_61 <= w_data;
        end
        if(_zz_2[62]) begin
          shift_q_map_62 <= w_data;
        end
        if(_zz_2[63]) begin
          shift_q_map_63 <= w_data;
        end
      end
    end
  end


endmodule

//MIMOReceiverUnit replaced by MIMOReceiverUnit

//MIMOReceiverUnit replaced by MIMOReceiverUnit

//MIMOReceiverUnit replaced by MIMOReceiverUnit

//MIMOReceiverUnit replaced by MIMOReceiverUnit

//MIMOReceiverUnit replaced by MIMOReceiverUnit

//MIMOReceiverUnit replaced by MIMOReceiverUnit

//MIMOReceiverUnit replaced by MIMOReceiverUnit

module MIMOReceiverUnit (
  input      [15:0]   shift_i_0,
  input      [15:0]   shift_i_1,
  input      [15:0]   shift_i_2,
  input      [15:0]   shift_i_3,
  input      [15:0]   shift_i_4,
  input      [15:0]   shift_i_5,
  input      [15:0]   shift_i_6,
  input      [15:0]   shift_i_7,
  input      [15:0]   shift_q_0,
  input      [15:0]   shift_q_1,
  input      [15:0]   shift_q_2,
  input      [15:0]   shift_q_3,
  input      [15:0]   shift_q_4,
  input      [15:0]   shift_q_5,
  input      [15:0]   shift_q_6,
  input      [15:0]   shift_q_7,
  input               mod_iq_valid,
  input      [15:0]   mod_iq_payload_cha_i,
  input      [15:0]   mod_iq_payload_cha_q,
  output              base_sub_iq_valid,
  output     [31:0]   base_sub_iq_payload_cha_i,
  output     [31:0]   base_sub_iq_payload_cha_q,
  input               rf_clk,
  input               rf_resetn
);

  wire       [31:0]   _zz_trans_i_vec_0;
  wire       [31:0]   _zz_trans_i_vec_0_1;
  wire       [31:0]   _zz_trans_q_vec_0;
  wire       [31:0]   _zz_trans_q_vec_0_1;
  wire       [31:0]   _zz_trans_i_vec_1;
  wire       [31:0]   _zz_trans_i_vec_1_1;
  wire       [31:0]   _zz_trans_q_vec_1;
  wire       [31:0]   _zz_trans_q_vec_1_1;
  wire       [31:0]   _zz_trans_i_vec_2;
  wire       [31:0]   _zz_trans_i_vec_2_1;
  wire       [31:0]   _zz_trans_q_vec_2;
  wire       [31:0]   _zz_trans_q_vec_2_1;
  wire       [31:0]   _zz_trans_i_vec_3;
  wire       [31:0]   _zz_trans_i_vec_3_1;
  wire       [31:0]   _zz_trans_q_vec_3;
  wire       [31:0]   _zz_trans_q_vec_3_1;
  wire       [31:0]   _zz_trans_i_vec_4;
  wire       [31:0]   _zz_trans_i_vec_4_1;
  wire       [31:0]   _zz_trans_q_vec_4;
  wire       [31:0]   _zz_trans_q_vec_4_1;
  wire       [31:0]   _zz_trans_i_vec_5;
  wire       [31:0]   _zz_trans_i_vec_5_1;
  wire       [31:0]   _zz_trans_q_vec_5;
  wire       [31:0]   _zz_trans_q_vec_5_1;
  wire       [31:0]   _zz_trans_i_vec_6;
  wire       [31:0]   _zz_trans_i_vec_6_1;
  wire       [31:0]   _zz_trans_q_vec_6;
  wire       [31:0]   _zz_trans_q_vec_6_1;
  wire       [31:0]   _zz_trans_i_vec_7;
  wire       [31:0]   _zz_trans_i_vec_7_1;
  wire       [31:0]   _zz_trans_q_vec_7;
  wire       [31:0]   _zz_trans_q_vec_7_1;
  wire       [30:0]   _zz__zz_base_sub_iq_payload_cha_i;
  wire       [31:0]   _zz__zz_base_sub_iq_payload_cha_i_1;
  wire       [30:0]   _zz__zz_base_sub_iq_payload_cha_i_1_1;
  wire       [31:0]   _zz__zz_base_sub_iq_payload_cha_i_1_2;
  wire       [30:0]   _zz__zz_base_sub_iq_payload_cha_i_2;
  wire       [31:0]   _zz__zz_base_sub_iq_payload_cha_i_2_1;
  wire       [30:0]   _zz__zz_base_sub_iq_payload_cha_i_3;
  wire       [31:0]   _zz__zz_base_sub_iq_payload_cha_i_3_1;
  wire       [30:0]   _zz__zz_base_sub_iq_payload_cha_i_4;
  wire       [31:0]   _zz__zz_base_sub_iq_payload_cha_i_4_1;
  wire       [30:0]   _zz__zz_base_sub_iq_payload_cha_i_5;
  wire       [31:0]   _zz__zz_base_sub_iq_payload_cha_i_5_1;
  wire       [30:0]   _zz__zz_base_sub_iq_payload_cha_i_6;
  wire       [31:0]   _zz__zz_base_sub_iq_payload_cha_i_6_1;
  wire       [30:0]   _zz__zz_base_sub_iq_payload_cha_q;
  wire       [31:0]   _zz__zz_base_sub_iq_payload_cha_q_1;
  wire       [30:0]   _zz__zz_base_sub_iq_payload_cha_q_1_1;
  wire       [31:0]   _zz__zz_base_sub_iq_payload_cha_q_1_2;
  wire       [30:0]   _zz__zz_base_sub_iq_payload_cha_q_2;
  wire       [31:0]   _zz__zz_base_sub_iq_payload_cha_q_2_1;
  wire       [30:0]   _zz__zz_base_sub_iq_payload_cha_q_3;
  wire       [31:0]   _zz__zz_base_sub_iq_payload_cha_q_3_1;
  wire       [30:0]   _zz__zz_base_sub_iq_payload_cha_q_4;
  wire       [31:0]   _zz__zz_base_sub_iq_payload_cha_q_4_1;
  wire       [30:0]   _zz__zz_base_sub_iq_payload_cha_q_5;
  wire       [31:0]   _zz__zz_base_sub_iq_payload_cha_q_5_1;
  wire       [30:0]   _zz__zz_base_sub_iq_payload_cha_q_6;
  wire       [31:0]   _zz__zz_base_sub_iq_payload_cha_q_6_1;
  reg        [15:0]   mod_iq_buf_cha_i;
  reg        [15:0]   mod_iq_buf_cha_q;
  reg                 mod_valid_buf;
  reg        [31:0]   trans_i_vec_0;
  reg        [31:0]   trans_i_vec_1;
  reg        [31:0]   trans_i_vec_2;
  reg        [31:0]   trans_i_vec_3;
  reg        [31:0]   trans_i_vec_4;
  reg        [31:0]   trans_i_vec_5;
  reg        [31:0]   trans_i_vec_6;
  reg        [31:0]   trans_i_vec_7;
  reg        [31:0]   trans_q_vec_0;
  reg        [31:0]   trans_q_vec_1;
  reg        [31:0]   trans_q_vec_2;
  reg        [31:0]   trans_q_vec_3;
  reg        [31:0]   trans_q_vec_4;
  reg        [31:0]   trans_q_vec_5;
  reg        [31:0]   trans_q_vec_6;
  reg        [31:0]   trans_q_vec_7;
  reg                 trans_valid;
  reg        [31:0]   _zz_base_sub_iq_payload_cha_i;
  reg        [31:0]   _zz_base_sub_iq_payload_cha_i_1;
  reg        [31:0]   _zz_base_sub_iq_payload_cha_i_2;
  reg        [31:0]   _zz_base_sub_iq_payload_cha_i_3;
  reg        [31:0]   _zz_base_sub_iq_payload_cha_i_4;
  reg        [31:0]   _zz_base_sub_iq_payload_cha_i_5;
  reg        [31:0]   _zz_base_sub_iq_payload_cha_i_6;
  reg        [31:0]   _zz_base_sub_iq_payload_cha_q;
  reg        [31:0]   _zz_base_sub_iq_payload_cha_q_1;
  reg        [31:0]   _zz_base_sub_iq_payload_cha_q_2;
  reg        [31:0]   _zz_base_sub_iq_payload_cha_q_3;
  reg        [31:0]   _zz_base_sub_iq_payload_cha_q_4;
  reg        [31:0]   _zz_base_sub_iq_payload_cha_q_5;
  reg        [31:0]   _zz_base_sub_iq_payload_cha_q_6;
  reg                 trans_valid_delay_1;
  reg                 trans_valid_delay_2;
  reg                 trans_valid_delay_3;

  assign _zz_trans_i_vec_0 = ($signed(mod_iq_buf_cha_i) * $signed(shift_i_0));
  assign _zz_trans_i_vec_0_1 = ($signed(mod_iq_buf_cha_q) * $signed(shift_q_0));
  assign _zz_trans_q_vec_0 = ($signed(mod_iq_buf_cha_i) * $signed(shift_q_0));
  assign _zz_trans_q_vec_0_1 = ($signed(mod_iq_buf_cha_q) * $signed(shift_i_0));
  assign _zz_trans_i_vec_1 = ($signed(mod_iq_buf_cha_i) * $signed(shift_i_1));
  assign _zz_trans_i_vec_1_1 = ($signed(mod_iq_buf_cha_q) * $signed(shift_q_1));
  assign _zz_trans_q_vec_1 = ($signed(mod_iq_buf_cha_i) * $signed(shift_q_1));
  assign _zz_trans_q_vec_1_1 = ($signed(mod_iq_buf_cha_q) * $signed(shift_i_1));
  assign _zz_trans_i_vec_2 = ($signed(mod_iq_buf_cha_i) * $signed(shift_i_2));
  assign _zz_trans_i_vec_2_1 = ($signed(mod_iq_buf_cha_q) * $signed(shift_q_2));
  assign _zz_trans_q_vec_2 = ($signed(mod_iq_buf_cha_i) * $signed(shift_q_2));
  assign _zz_trans_q_vec_2_1 = ($signed(mod_iq_buf_cha_q) * $signed(shift_i_2));
  assign _zz_trans_i_vec_3 = ($signed(mod_iq_buf_cha_i) * $signed(shift_i_3));
  assign _zz_trans_i_vec_3_1 = ($signed(mod_iq_buf_cha_q) * $signed(shift_q_3));
  assign _zz_trans_q_vec_3 = ($signed(mod_iq_buf_cha_i) * $signed(shift_q_3));
  assign _zz_trans_q_vec_3_1 = ($signed(mod_iq_buf_cha_q) * $signed(shift_i_3));
  assign _zz_trans_i_vec_4 = ($signed(mod_iq_buf_cha_i) * $signed(shift_i_4));
  assign _zz_trans_i_vec_4_1 = ($signed(mod_iq_buf_cha_q) * $signed(shift_q_4));
  assign _zz_trans_q_vec_4 = ($signed(mod_iq_buf_cha_i) * $signed(shift_q_4));
  assign _zz_trans_q_vec_4_1 = ($signed(mod_iq_buf_cha_q) * $signed(shift_i_4));
  assign _zz_trans_i_vec_5 = ($signed(mod_iq_buf_cha_i) * $signed(shift_i_5));
  assign _zz_trans_i_vec_5_1 = ($signed(mod_iq_buf_cha_q) * $signed(shift_q_5));
  assign _zz_trans_q_vec_5 = ($signed(mod_iq_buf_cha_i) * $signed(shift_q_5));
  assign _zz_trans_q_vec_5_1 = ($signed(mod_iq_buf_cha_q) * $signed(shift_i_5));
  assign _zz_trans_i_vec_6 = ($signed(mod_iq_buf_cha_i) * $signed(shift_i_6));
  assign _zz_trans_i_vec_6_1 = ($signed(mod_iq_buf_cha_q) * $signed(shift_q_6));
  assign _zz_trans_q_vec_6 = ($signed(mod_iq_buf_cha_i) * $signed(shift_q_6));
  assign _zz_trans_q_vec_6_1 = ($signed(mod_iq_buf_cha_q) * $signed(shift_i_6));
  assign _zz_trans_i_vec_7 = ($signed(mod_iq_buf_cha_i) * $signed(shift_i_7));
  assign _zz_trans_i_vec_7_1 = ($signed(mod_iq_buf_cha_q) * $signed(shift_q_7));
  assign _zz_trans_q_vec_7 = ($signed(mod_iq_buf_cha_i) * $signed(shift_q_7));
  assign _zz_trans_q_vec_7_1 = ($signed(mod_iq_buf_cha_q) * $signed(shift_i_7));
  assign _zz__zz_base_sub_iq_payload_cha_i = (_zz__zz_base_sub_iq_payload_cha_i_1 >>> 1);
  assign _zz__zz_base_sub_iq_payload_cha_i_1 = ($signed(trans_i_vec_0) + $signed(trans_i_vec_1));
  assign _zz__zz_base_sub_iq_payload_cha_i_1_1 = (_zz__zz_base_sub_iq_payload_cha_i_1_2 >>> 1);
  assign _zz__zz_base_sub_iq_payload_cha_i_1_2 = ($signed(trans_i_vec_2) + $signed(trans_i_vec_3));
  assign _zz__zz_base_sub_iq_payload_cha_i_2 = (_zz__zz_base_sub_iq_payload_cha_i_2_1 >>> 1);
  assign _zz__zz_base_sub_iq_payload_cha_i_2_1 = ($signed(trans_i_vec_4) + $signed(trans_i_vec_5));
  assign _zz__zz_base_sub_iq_payload_cha_i_3 = (_zz__zz_base_sub_iq_payload_cha_i_3_1 >>> 1);
  assign _zz__zz_base_sub_iq_payload_cha_i_3_1 = ($signed(trans_i_vec_6) + $signed(trans_i_vec_7));
  assign _zz__zz_base_sub_iq_payload_cha_i_4 = (_zz__zz_base_sub_iq_payload_cha_i_4_1 >>> 1);
  assign _zz__zz_base_sub_iq_payload_cha_i_4_1 = ($signed(_zz_base_sub_iq_payload_cha_i) + $signed(_zz_base_sub_iq_payload_cha_i_1));
  assign _zz__zz_base_sub_iq_payload_cha_i_5 = (_zz__zz_base_sub_iq_payload_cha_i_5_1 >>> 1);
  assign _zz__zz_base_sub_iq_payload_cha_i_5_1 = ($signed(_zz_base_sub_iq_payload_cha_i_2) + $signed(_zz_base_sub_iq_payload_cha_i_3));
  assign _zz__zz_base_sub_iq_payload_cha_i_6 = (_zz__zz_base_sub_iq_payload_cha_i_6_1 >>> 1);
  assign _zz__zz_base_sub_iq_payload_cha_i_6_1 = ($signed(_zz_base_sub_iq_payload_cha_i_4) + $signed(_zz_base_sub_iq_payload_cha_i_5));
  assign _zz__zz_base_sub_iq_payload_cha_q = (_zz__zz_base_sub_iq_payload_cha_q_1 >>> 1);
  assign _zz__zz_base_sub_iq_payload_cha_q_1 = ($signed(trans_q_vec_0) + $signed(trans_q_vec_1));
  assign _zz__zz_base_sub_iq_payload_cha_q_1_1 = (_zz__zz_base_sub_iq_payload_cha_q_1_2 >>> 1);
  assign _zz__zz_base_sub_iq_payload_cha_q_1_2 = ($signed(trans_q_vec_2) + $signed(trans_q_vec_3));
  assign _zz__zz_base_sub_iq_payload_cha_q_2 = (_zz__zz_base_sub_iq_payload_cha_q_2_1 >>> 1);
  assign _zz__zz_base_sub_iq_payload_cha_q_2_1 = ($signed(trans_q_vec_4) + $signed(trans_q_vec_5));
  assign _zz__zz_base_sub_iq_payload_cha_q_3 = (_zz__zz_base_sub_iq_payload_cha_q_3_1 >>> 1);
  assign _zz__zz_base_sub_iq_payload_cha_q_3_1 = ($signed(trans_q_vec_6) + $signed(trans_q_vec_7));
  assign _zz__zz_base_sub_iq_payload_cha_q_4 = (_zz__zz_base_sub_iq_payload_cha_q_4_1 >>> 1);
  assign _zz__zz_base_sub_iq_payload_cha_q_4_1 = ($signed(_zz_base_sub_iq_payload_cha_q) + $signed(_zz_base_sub_iq_payload_cha_q_1));
  assign _zz__zz_base_sub_iq_payload_cha_q_5 = (_zz__zz_base_sub_iq_payload_cha_q_5_1 >>> 1);
  assign _zz__zz_base_sub_iq_payload_cha_q_5_1 = ($signed(_zz_base_sub_iq_payload_cha_q_2) + $signed(_zz_base_sub_iq_payload_cha_q_3));
  assign _zz__zz_base_sub_iq_payload_cha_q_6 = (_zz__zz_base_sub_iq_payload_cha_q_6_1 >>> 1);
  assign _zz__zz_base_sub_iq_payload_cha_q_6_1 = ($signed(_zz_base_sub_iq_payload_cha_q_4) + $signed(_zz_base_sub_iq_payload_cha_q_5));
  assign base_sub_iq_payload_cha_i = _zz_base_sub_iq_payload_cha_i_6;
  assign base_sub_iq_payload_cha_q = _zz_base_sub_iq_payload_cha_q_6;
  assign base_sub_iq_valid = trans_valid_delay_3;
  always @(posedge rf_clk) begin
    mod_iq_buf_cha_i <= mod_iq_payload_cha_i;
    mod_iq_buf_cha_q <= mod_iq_payload_cha_q;
    if(mod_valid_buf) begin
      trans_i_vec_0 <= ($signed(_zz_trans_i_vec_0) - $signed(_zz_trans_i_vec_0_1));
      trans_q_vec_0 <= ($signed(_zz_trans_q_vec_0) + $signed(_zz_trans_q_vec_0_1));
      trans_i_vec_1 <= ($signed(_zz_trans_i_vec_1) - $signed(_zz_trans_i_vec_1_1));
      trans_q_vec_1 <= ($signed(_zz_trans_q_vec_1) + $signed(_zz_trans_q_vec_1_1));
      trans_i_vec_2 <= ($signed(_zz_trans_i_vec_2) - $signed(_zz_trans_i_vec_2_1));
      trans_q_vec_2 <= ($signed(_zz_trans_q_vec_2) + $signed(_zz_trans_q_vec_2_1));
      trans_i_vec_3 <= ($signed(_zz_trans_i_vec_3) - $signed(_zz_trans_i_vec_3_1));
      trans_q_vec_3 <= ($signed(_zz_trans_q_vec_3) + $signed(_zz_trans_q_vec_3_1));
      trans_i_vec_4 <= ($signed(_zz_trans_i_vec_4) - $signed(_zz_trans_i_vec_4_1));
      trans_q_vec_4 <= ($signed(_zz_trans_q_vec_4) + $signed(_zz_trans_q_vec_4_1));
      trans_i_vec_5 <= ($signed(_zz_trans_i_vec_5) - $signed(_zz_trans_i_vec_5_1));
      trans_q_vec_5 <= ($signed(_zz_trans_q_vec_5) + $signed(_zz_trans_q_vec_5_1));
      trans_i_vec_6 <= ($signed(_zz_trans_i_vec_6) - $signed(_zz_trans_i_vec_6_1));
      trans_q_vec_6 <= ($signed(_zz_trans_q_vec_6) + $signed(_zz_trans_q_vec_6_1));
      trans_i_vec_7 <= ($signed(_zz_trans_i_vec_7) - $signed(_zz_trans_i_vec_7_1));
      trans_q_vec_7 <= ($signed(_zz_trans_q_vec_7) + $signed(_zz_trans_q_vec_7_1));
    end else begin
      trans_i_vec_0 <= 32'h0;
      trans_q_vec_0 <= 32'h0;
      trans_i_vec_1 <= 32'h0;
      trans_q_vec_1 <= 32'h0;
      trans_i_vec_2 <= 32'h0;
      trans_q_vec_2 <= 32'h0;
      trans_i_vec_3 <= 32'h0;
      trans_q_vec_3 <= 32'h0;
      trans_i_vec_4 <= 32'h0;
      trans_q_vec_4 <= 32'h0;
      trans_i_vec_5 <= 32'h0;
      trans_q_vec_5 <= 32'h0;
      trans_i_vec_6 <= 32'h0;
      trans_q_vec_6 <= 32'h0;
      trans_i_vec_7 <= 32'h0;
      trans_q_vec_7 <= 32'h0;
    end
    _zz_base_sub_iq_payload_cha_i <= {{1{_zz__zz_base_sub_iq_payload_cha_i[30]}}, _zz__zz_base_sub_iq_payload_cha_i};
    _zz_base_sub_iq_payload_cha_i_1 <= {{1{_zz__zz_base_sub_iq_payload_cha_i_1_1[30]}}, _zz__zz_base_sub_iq_payload_cha_i_1_1};
    _zz_base_sub_iq_payload_cha_i_2 <= {{1{_zz__zz_base_sub_iq_payload_cha_i_2[30]}}, _zz__zz_base_sub_iq_payload_cha_i_2};
    _zz_base_sub_iq_payload_cha_i_3 <= {{1{_zz__zz_base_sub_iq_payload_cha_i_3[30]}}, _zz__zz_base_sub_iq_payload_cha_i_3};
    _zz_base_sub_iq_payload_cha_i_4 <= {{1{_zz__zz_base_sub_iq_payload_cha_i_4[30]}}, _zz__zz_base_sub_iq_payload_cha_i_4};
    _zz_base_sub_iq_payload_cha_i_5 <= {{1{_zz__zz_base_sub_iq_payload_cha_i_5[30]}}, _zz__zz_base_sub_iq_payload_cha_i_5};
    _zz_base_sub_iq_payload_cha_i_6 <= {{1{_zz__zz_base_sub_iq_payload_cha_i_6[30]}}, _zz__zz_base_sub_iq_payload_cha_i_6};
    _zz_base_sub_iq_payload_cha_q <= {{1{_zz__zz_base_sub_iq_payload_cha_q[30]}}, _zz__zz_base_sub_iq_payload_cha_q};
    _zz_base_sub_iq_payload_cha_q_1 <= {{1{_zz__zz_base_sub_iq_payload_cha_q_1_1[30]}}, _zz__zz_base_sub_iq_payload_cha_q_1_1};
    _zz_base_sub_iq_payload_cha_q_2 <= {{1{_zz__zz_base_sub_iq_payload_cha_q_2[30]}}, _zz__zz_base_sub_iq_payload_cha_q_2};
    _zz_base_sub_iq_payload_cha_q_3 <= {{1{_zz__zz_base_sub_iq_payload_cha_q_3[30]}}, _zz__zz_base_sub_iq_payload_cha_q_3};
    _zz_base_sub_iq_payload_cha_q_4 <= {{1{_zz__zz_base_sub_iq_payload_cha_q_4[30]}}, _zz__zz_base_sub_iq_payload_cha_q_4};
    _zz_base_sub_iq_payload_cha_q_5 <= {{1{_zz__zz_base_sub_iq_payload_cha_q_5[30]}}, _zz__zz_base_sub_iq_payload_cha_q_5};
    _zz_base_sub_iq_payload_cha_q_6 <= {{1{_zz__zz_base_sub_iq_payload_cha_q_6[30]}}, _zz__zz_base_sub_iq_payload_cha_q_6};
    trans_valid_delay_1 <= trans_valid;
    trans_valid_delay_2 <= trans_valid_delay_1;
    trans_valid_delay_3 <= trans_valid_delay_2;
  end

  always @(posedge rf_clk) begin
    if(!rf_resetn) begin
      mod_valid_buf <= 1'b0;
      trans_valid <= 1'b0;
    end else begin
      mod_valid_buf <= mod_iq_valid;
      if(mod_valid_buf) begin
        trans_valid <= 1'b1;
      end else begin
        trans_valid <= 1'b0;
      end
    end
  end


endmodule
