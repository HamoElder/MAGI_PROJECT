// Generator : SpinalHDL v1.6.0    git head : 73c8d8e2b86b45646e9d0b2e729291f2b65e6be3
// Component : UnsignedDivider
// Git hash  : 090aef073dde5541acfdebf275d47dcc675b45b6



module UnsignedDivider (
  input               flush,
  input               cmd_valid,
  output              cmd_ready,
  input      [15:0]   cmd_payload_numerator,
  input      [15:0]   cmd_payload_denominator,
  output              rsp_valid,
  input               rsp_ready,
  output     [15:0]   rsp_payload_quotient,
  output     [15:0]   rsp_payload_remainder,
  output              rsp_payload_error,
  input               clk,
  input               reset
);
  wire       [16:0]   _zz__zz_rsp_payload_quotient_61;
  wire       [16:0]   _zz__zz_rsp_payload_quotient_62;
  wire       [16:0]   _zz__zz_rsp_payload_quotient_63;
  wire       [16:0]   _zz__zz_rsp_payload_quotient_64;
  wire       [16:0]   _zz__zz_rsp_payload_quotient_65;
  wire       [16:0]   _zz__zz_rsp_payload_quotient_66;
  wire       [16:0]   _zz__zz_rsp_payload_quotient_67;
  wire       [16:0]   _zz__zz_rsp_payload_quotient_68;
  wire       [16:0]   _zz__zz_rsp_payload_quotient_69;
  wire       [16:0]   _zz__zz_rsp_payload_quotient_70;
  wire       [16:0]   _zz__zz_rsp_payload_quotient_71;
  wire       [16:0]   _zz__zz_rsp_payload_quotient_72;
  wire       [16:0]   _zz__zz_rsp_payload_quotient_73;
  wire       [16:0]   _zz__zz_rsp_payload_quotient_74;
  wire       [16:0]   _zz__zz_rsp_payload_quotient_75;
  wire       [16:0]   _zz__zz_rsp_payload_quotient_1;
  wire       [16:0]   _zz__zz_rsp_payload_quotient_2;
  wire       [16:0]   _zz__zz_rsp_payload_quotient_3;
  wire       [16:0]   _zz__zz_rsp_payload_quotient_4;
  wire       [16:0]   _zz__zz_rsp_payload_quotient_5;
  wire       [16:0]   _zz__zz_rsp_payload_quotient_6;
  wire       [16:0]   _zz__zz_rsp_payload_quotient_7;
  wire       [16:0]   _zz__zz_rsp_payload_quotient_8;
  wire       [16:0]   _zz__zz_rsp_payload_quotient_9;
  wire       [16:0]   _zz__zz_rsp_payload_quotient_10;
  wire       [16:0]   _zz__zz_rsp_payload_quotient_11;
  wire       [16:0]   _zz__zz_rsp_payload_quotient_12;
  wire       [16:0]   _zz__zz_rsp_payload_quotient_13;
  wire       [16:0]   _zz__zz_rsp_payload_quotient_14;
  wire       [16:0]   _zz__zz_rsp_payload_quotient_15;
  reg                 _zz_rsp_valid;
  reg                 _zz_rsp_valid_1;
  reg                 _zz_rsp_valid_2;
  reg                 _zz_rsp_valid_3;
  reg                 _zz_rsp_valid_4;
  reg                 _zz_rsp_valid_5;
  reg                 _zz_rsp_valid_6;
  reg                 _zz_rsp_valid_7;
  reg                 _zz_rsp_valid_8;
  reg                 _zz_rsp_valid_9;
  reg                 _zz_rsp_valid_10;
  reg                 _zz_rsp_valid_11;
  reg                 _zz_rsp_valid_12;
  reg                 _zz_rsp_valid_13;
  reg                 _zz_rsp_valid_14;
  reg                 _zz_rsp_valid_15;
  reg        [15:0]   _zz_rsp_payload_quotient;
  reg        [15:0]   _zz_rsp_payload_quotient_1;
  reg        [15:0]   _zz_rsp_payload_quotient_2;
  reg        [15:0]   _zz_rsp_payload_quotient_3;
  reg        [15:0]   _zz_rsp_payload_quotient_4;
  reg        [15:0]   _zz_rsp_payload_quotient_5;
  reg        [15:0]   _zz_rsp_payload_quotient_6;
  reg        [15:0]   _zz_rsp_payload_quotient_7;
  reg        [15:0]   _zz_rsp_payload_quotient_8;
  reg        [15:0]   _zz_rsp_payload_quotient_9;
  reg        [15:0]   _zz_rsp_payload_quotient_10;
  reg        [15:0]   _zz_rsp_payload_quotient_11;
  reg        [15:0]   _zz_rsp_payload_quotient_12;
  reg        [15:0]   _zz_rsp_payload_quotient_13;
  reg        [15:0]   _zz_rsp_payload_quotient_14;
  reg        [15:0]   _zz_rsp_payload_quotient_15;
  reg        [15:0]   _zz_rsp_payload_quotient_16;
  reg        [15:0]   _zz_rsp_payload_quotient_17;
  reg        [15:0]   _zz_rsp_payload_quotient_18;
  reg        [15:0]   _zz_rsp_payload_quotient_19;
  reg        [15:0]   _zz_rsp_payload_quotient_20;
  reg        [15:0]   _zz_rsp_payload_quotient_21;
  reg        [15:0]   _zz_rsp_payload_quotient_22;
  reg        [15:0]   _zz_rsp_payload_quotient_23;
  reg        [15:0]   _zz_rsp_payload_quotient_24;
  reg        [15:0]   _zz_rsp_payload_quotient_25;
  reg        [15:0]   _zz_rsp_payload_quotient_26;
  reg        [15:0]   _zz_rsp_payload_quotient_27;
  reg        [15:0]   _zz_rsp_payload_quotient_28;
  reg        [15:0]   _zz_rsp_payload_quotient_29;
  reg        [15:0]   _zz_rsp_payload_quotient_30;
  reg        [15:0]   _zz_rsp_payload_error;
  reg        [15:0]   _zz_rsp_payload_quotient_31;
  reg        [15:0]   _zz_rsp_payload_quotient_32;
  reg        [15:0]   _zz_rsp_payload_quotient_33;
  reg        [15:0]   _zz_rsp_payload_quotient_34;
  reg        [15:0]   _zz_rsp_payload_quotient_35;
  reg        [15:0]   _zz_rsp_payload_quotient_36;
  reg        [15:0]   _zz_rsp_payload_quotient_37;
  reg        [15:0]   _zz_rsp_payload_quotient_38;
  reg        [15:0]   _zz_rsp_payload_quotient_39;
  reg        [15:0]   _zz_rsp_payload_quotient_40;
  reg        [15:0]   _zz_rsp_payload_quotient_41;
  reg        [15:0]   _zz_rsp_payload_quotient_42;
  reg        [15:0]   _zz_rsp_payload_quotient_43;
  reg        [15:0]   _zz_rsp_payload_quotient_44;
  reg        [15:0]   _zz_rsp_payload_quotient_45;
  reg        [15:0]   _zz_rsp_payload_remainder;
  wire       [16:0]   _zz_rsp_payload_quotient_46;
  wire       [16:0]   _zz_rsp_payload_quotient_47;
  wire       [16:0]   _zz_rsp_payload_quotient_48;
  wire       [16:0]   _zz_rsp_payload_quotient_49;
  wire       [16:0]   _zz_rsp_payload_quotient_50;
  wire       [16:0]   _zz_rsp_payload_quotient_51;
  wire       [16:0]   _zz_rsp_payload_quotient_52;
  wire       [16:0]   _zz_rsp_payload_quotient_53;
  wire       [16:0]   _zz_rsp_payload_quotient_54;
  wire       [16:0]   _zz_rsp_payload_quotient_55;
  wire       [16:0]   _zz_rsp_payload_quotient_56;
  wire       [16:0]   _zz_rsp_payload_quotient_57;
  wire       [16:0]   _zz_rsp_payload_quotient_58;
  wire       [16:0]   _zz_rsp_payload_quotient_59;
  wire       [16:0]   _zz_rsp_payload_quotient_60;
  wire       [16:0]   _zz_rsp_payload_quotient_61;
  wire       [16:0]   _zz_rsp_payload_quotient_62;
  wire       [16:0]   _zz_rsp_payload_quotient_63;
  wire       [16:0]   _zz_rsp_payload_quotient_64;
  wire       [16:0]   _zz_rsp_payload_quotient_65;
  wire       [16:0]   _zz_rsp_payload_quotient_66;
  wire       [16:0]   _zz_rsp_payload_quotient_67;
  wire       [16:0]   _zz_rsp_payload_quotient_68;
  wire       [16:0]   _zz_rsp_payload_quotient_69;
  wire       [16:0]   _zz_rsp_payload_quotient_70;
  wire       [16:0]   _zz_rsp_payload_quotient_71;
  wire       [16:0]   _zz_rsp_payload_quotient_72;
  wire       [16:0]   _zz_rsp_payload_quotient_73;
  wire       [16:0]   _zz_rsp_payload_quotient_74;
  wire       [16:0]   _zz_rsp_payload_quotient_75;
  wire                cmd_fire;
  wire                when_UnsignedDivider_l58;
  wire                when_UnsignedDivider_l58_1;
  wire                when_UnsignedDivider_l58_2;
  wire                when_UnsignedDivider_l58_3;
  wire                when_UnsignedDivider_l58_4;
  wire                when_UnsignedDivider_l58_5;
  wire                when_UnsignedDivider_l58_6;
  wire                when_UnsignedDivider_l58_7;
  wire                when_UnsignedDivider_l58_8;
  wire                when_UnsignedDivider_l58_9;
  wire                when_UnsignedDivider_l58_10;
  wire                when_UnsignedDivider_l58_11;
  wire                when_UnsignedDivider_l58_12;
  wire                when_UnsignedDivider_l58_13;
  wire                when_UnsignedDivider_l58_14;

  assign _zz__zz_rsp_payload_quotient_61 = {1'd0, _zz_rsp_payload_quotient_16};
  assign _zz__zz_rsp_payload_quotient_62 = {1'd0, _zz_rsp_payload_quotient_17};
  assign _zz__zz_rsp_payload_quotient_63 = {1'd0, _zz_rsp_payload_quotient_18};
  assign _zz__zz_rsp_payload_quotient_64 = {1'd0, _zz_rsp_payload_quotient_19};
  assign _zz__zz_rsp_payload_quotient_65 = {1'd0, _zz_rsp_payload_quotient_20};
  assign _zz__zz_rsp_payload_quotient_66 = {1'd0, _zz_rsp_payload_quotient_21};
  assign _zz__zz_rsp_payload_quotient_67 = {1'd0, _zz_rsp_payload_quotient_22};
  assign _zz__zz_rsp_payload_quotient_68 = {1'd0, _zz_rsp_payload_quotient_23};
  assign _zz__zz_rsp_payload_quotient_69 = {1'd0, _zz_rsp_payload_quotient_24};
  assign _zz__zz_rsp_payload_quotient_70 = {1'd0, _zz_rsp_payload_quotient_25};
  assign _zz__zz_rsp_payload_quotient_71 = {1'd0, _zz_rsp_payload_quotient_26};
  assign _zz__zz_rsp_payload_quotient_72 = {1'd0, _zz_rsp_payload_quotient_27};
  assign _zz__zz_rsp_payload_quotient_73 = {1'd0, _zz_rsp_payload_quotient_28};
  assign _zz__zz_rsp_payload_quotient_74 = {1'd0, _zz_rsp_payload_quotient_29};
  assign _zz__zz_rsp_payload_quotient_75 = {1'd0, _zz_rsp_payload_quotient_30};
  assign _zz__zz_rsp_payload_quotient_1 = {_zz_rsp_payload_quotient,(! _zz_rsp_payload_quotient_61[16])};
  assign _zz__zz_rsp_payload_quotient_2 = {_zz_rsp_payload_quotient_1,(! _zz_rsp_payload_quotient_62[16])};
  assign _zz__zz_rsp_payload_quotient_3 = {_zz_rsp_payload_quotient_2,(! _zz_rsp_payload_quotient_63[16])};
  assign _zz__zz_rsp_payload_quotient_4 = {_zz_rsp_payload_quotient_3,(! _zz_rsp_payload_quotient_64[16])};
  assign _zz__zz_rsp_payload_quotient_5 = {_zz_rsp_payload_quotient_4,(! _zz_rsp_payload_quotient_65[16])};
  assign _zz__zz_rsp_payload_quotient_6 = {_zz_rsp_payload_quotient_5,(! _zz_rsp_payload_quotient_66[16])};
  assign _zz__zz_rsp_payload_quotient_7 = {_zz_rsp_payload_quotient_6,(! _zz_rsp_payload_quotient_67[16])};
  assign _zz__zz_rsp_payload_quotient_8 = {_zz_rsp_payload_quotient_7,(! _zz_rsp_payload_quotient_68[16])};
  assign _zz__zz_rsp_payload_quotient_9 = {_zz_rsp_payload_quotient_8,(! _zz_rsp_payload_quotient_69[16])};
  assign _zz__zz_rsp_payload_quotient_10 = {_zz_rsp_payload_quotient_9,(! _zz_rsp_payload_quotient_70[16])};
  assign _zz__zz_rsp_payload_quotient_11 = {_zz_rsp_payload_quotient_10,(! _zz_rsp_payload_quotient_71[16])};
  assign _zz__zz_rsp_payload_quotient_12 = {_zz_rsp_payload_quotient_11,(! _zz_rsp_payload_quotient_72[16])};
  assign _zz__zz_rsp_payload_quotient_13 = {_zz_rsp_payload_quotient_12,(! _zz_rsp_payload_quotient_73[16])};
  assign _zz__zz_rsp_payload_quotient_14 = {_zz_rsp_payload_quotient_13,(! _zz_rsp_payload_quotient_74[16])};
  assign _zz__zz_rsp_payload_quotient_15 = {_zz_rsp_payload_quotient_14,(! _zz_rsp_payload_quotient_75[16])};
  assign _zz_rsp_payload_quotient_46 = {_zz_rsp_payload_quotient_31,_zz_rsp_payload_quotient[15]};
  assign _zz_rsp_payload_quotient_61 = (_zz_rsp_payload_quotient_46 - _zz__zz_rsp_payload_quotient_61);
  assign _zz_rsp_payload_quotient_47 = {_zz_rsp_payload_quotient_32,_zz_rsp_payload_quotient_1[15]};
  assign _zz_rsp_payload_quotient_62 = (_zz_rsp_payload_quotient_47 - _zz__zz_rsp_payload_quotient_62);
  assign _zz_rsp_payload_quotient_48 = {_zz_rsp_payload_quotient_33,_zz_rsp_payload_quotient_2[15]};
  assign _zz_rsp_payload_quotient_63 = (_zz_rsp_payload_quotient_48 - _zz__zz_rsp_payload_quotient_63);
  assign _zz_rsp_payload_quotient_49 = {_zz_rsp_payload_quotient_34,_zz_rsp_payload_quotient_3[15]};
  assign _zz_rsp_payload_quotient_64 = (_zz_rsp_payload_quotient_49 - _zz__zz_rsp_payload_quotient_64);
  assign _zz_rsp_payload_quotient_50 = {_zz_rsp_payload_quotient_35,_zz_rsp_payload_quotient_4[15]};
  assign _zz_rsp_payload_quotient_65 = (_zz_rsp_payload_quotient_50 - _zz__zz_rsp_payload_quotient_65);
  assign _zz_rsp_payload_quotient_51 = {_zz_rsp_payload_quotient_36,_zz_rsp_payload_quotient_5[15]};
  assign _zz_rsp_payload_quotient_66 = (_zz_rsp_payload_quotient_51 - _zz__zz_rsp_payload_quotient_66);
  assign _zz_rsp_payload_quotient_52 = {_zz_rsp_payload_quotient_37,_zz_rsp_payload_quotient_6[15]};
  assign _zz_rsp_payload_quotient_67 = (_zz_rsp_payload_quotient_52 - _zz__zz_rsp_payload_quotient_67);
  assign _zz_rsp_payload_quotient_53 = {_zz_rsp_payload_quotient_38,_zz_rsp_payload_quotient_7[15]};
  assign _zz_rsp_payload_quotient_68 = (_zz_rsp_payload_quotient_53 - _zz__zz_rsp_payload_quotient_68);
  assign _zz_rsp_payload_quotient_54 = {_zz_rsp_payload_quotient_39,_zz_rsp_payload_quotient_8[15]};
  assign _zz_rsp_payload_quotient_69 = (_zz_rsp_payload_quotient_54 - _zz__zz_rsp_payload_quotient_69);
  assign _zz_rsp_payload_quotient_55 = {_zz_rsp_payload_quotient_40,_zz_rsp_payload_quotient_9[15]};
  assign _zz_rsp_payload_quotient_70 = (_zz_rsp_payload_quotient_55 - _zz__zz_rsp_payload_quotient_70);
  assign _zz_rsp_payload_quotient_56 = {_zz_rsp_payload_quotient_41,_zz_rsp_payload_quotient_10[15]};
  assign _zz_rsp_payload_quotient_71 = (_zz_rsp_payload_quotient_56 - _zz__zz_rsp_payload_quotient_71);
  assign _zz_rsp_payload_quotient_57 = {_zz_rsp_payload_quotient_42,_zz_rsp_payload_quotient_11[15]};
  assign _zz_rsp_payload_quotient_72 = (_zz_rsp_payload_quotient_57 - _zz__zz_rsp_payload_quotient_72);
  assign _zz_rsp_payload_quotient_58 = {_zz_rsp_payload_quotient_43,_zz_rsp_payload_quotient_12[15]};
  assign _zz_rsp_payload_quotient_73 = (_zz_rsp_payload_quotient_58 - _zz__zz_rsp_payload_quotient_73);
  assign _zz_rsp_payload_quotient_59 = {_zz_rsp_payload_quotient_44,_zz_rsp_payload_quotient_13[15]};
  assign _zz_rsp_payload_quotient_74 = (_zz_rsp_payload_quotient_59 - _zz__zz_rsp_payload_quotient_74);
  assign _zz_rsp_payload_quotient_60 = {_zz_rsp_payload_quotient_45,_zz_rsp_payload_quotient_14[15]};
  assign _zz_rsp_payload_quotient_75 = (_zz_rsp_payload_quotient_60 - _zz__zz_rsp_payload_quotient_75);
  assign cmd_ready = rsp_ready;
  assign cmd_fire = (cmd_valid && cmd_ready);
  assign when_UnsignedDivider_l58 = (! _zz_rsp_payload_quotient_61[16]);
  assign when_UnsignedDivider_l58_1 = (! _zz_rsp_payload_quotient_62[16]);
  assign when_UnsignedDivider_l58_2 = (! _zz_rsp_payload_quotient_63[16]);
  assign when_UnsignedDivider_l58_3 = (! _zz_rsp_payload_quotient_64[16]);
  assign when_UnsignedDivider_l58_4 = (! _zz_rsp_payload_quotient_65[16]);
  assign when_UnsignedDivider_l58_5 = (! _zz_rsp_payload_quotient_66[16]);
  assign when_UnsignedDivider_l58_6 = (! _zz_rsp_payload_quotient_67[16]);
  assign when_UnsignedDivider_l58_7 = (! _zz_rsp_payload_quotient_68[16]);
  assign when_UnsignedDivider_l58_8 = (! _zz_rsp_payload_quotient_69[16]);
  assign when_UnsignedDivider_l58_9 = (! _zz_rsp_payload_quotient_70[16]);
  assign when_UnsignedDivider_l58_10 = (! _zz_rsp_payload_quotient_71[16]);
  assign when_UnsignedDivider_l58_11 = (! _zz_rsp_payload_quotient_72[16]);
  assign when_UnsignedDivider_l58_12 = (! _zz_rsp_payload_quotient_73[16]);
  assign when_UnsignedDivider_l58_13 = (! _zz_rsp_payload_quotient_74[16]);
  assign when_UnsignedDivider_l58_14 = (! _zz_rsp_payload_quotient_75[16]);
  assign rsp_valid = _zz_rsp_valid_15;
  assign rsp_payload_quotient = _zz_rsp_payload_quotient_15;
  assign rsp_payload_remainder = _zz_rsp_payload_remainder;
  assign rsp_payload_error = (_zz_rsp_payload_error == 16'h0);
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _zz_rsp_valid <= 1'b0;
      _zz_rsp_valid_1 <= 1'b0;
      _zz_rsp_valid_2 <= 1'b0;
      _zz_rsp_valid_3 <= 1'b0;
      _zz_rsp_valid_4 <= 1'b0;
      _zz_rsp_valid_5 <= 1'b0;
      _zz_rsp_valid_6 <= 1'b0;
      _zz_rsp_valid_7 <= 1'b0;
      _zz_rsp_valid_8 <= 1'b0;
      _zz_rsp_valid_9 <= 1'b0;
      _zz_rsp_valid_10 <= 1'b0;
      _zz_rsp_valid_11 <= 1'b0;
      _zz_rsp_valid_12 <= 1'b0;
      _zz_rsp_valid_13 <= 1'b0;
      _zz_rsp_valid_14 <= 1'b0;
      _zz_rsp_valid_15 <= 1'b0;
    end else begin
      _zz_rsp_valid <= (flush ? 1'b0 : cmd_fire);
      _zz_rsp_valid_1 <= (flush ? 1'b0 : _zz_rsp_valid);
      _zz_rsp_valid_2 <= (flush ? 1'b0 : _zz_rsp_valid_1);
      _zz_rsp_valid_3 <= (flush ? 1'b0 : _zz_rsp_valid_2);
      _zz_rsp_valid_4 <= (flush ? 1'b0 : _zz_rsp_valid_3);
      _zz_rsp_valid_5 <= (flush ? 1'b0 : _zz_rsp_valid_4);
      _zz_rsp_valid_6 <= (flush ? 1'b0 : _zz_rsp_valid_5);
      _zz_rsp_valid_7 <= (flush ? 1'b0 : _zz_rsp_valid_6);
      _zz_rsp_valid_8 <= (flush ? 1'b0 : _zz_rsp_valid_7);
      _zz_rsp_valid_9 <= (flush ? 1'b0 : _zz_rsp_valid_8);
      _zz_rsp_valid_10 <= (flush ? 1'b0 : _zz_rsp_valid_9);
      _zz_rsp_valid_11 <= (flush ? 1'b0 : _zz_rsp_valid_10);
      _zz_rsp_valid_12 <= (flush ? 1'b0 : _zz_rsp_valid_11);
      _zz_rsp_valid_13 <= (flush ? 1'b0 : _zz_rsp_valid_12);
      _zz_rsp_valid_14 <= (flush ? 1'b0 : _zz_rsp_valid_13);
      _zz_rsp_valid_15 <= (flush ? 1'b0 : _zz_rsp_valid_14);
    end
  end

  always @(posedge clk) begin
    _zz_rsp_payload_quotient_16 <= cmd_payload_denominator;
    _zz_rsp_payload_quotient_31 <= 16'h0;
    _zz_rsp_payload_quotient <= cmd_payload_numerator;
    _zz_rsp_payload_quotient_17 <= _zz_rsp_payload_quotient_16;
    _zz_rsp_payload_quotient_1 <= _zz__zz_rsp_payload_quotient_1[15:0];
    if(when_UnsignedDivider_l58) begin
      _zz_rsp_payload_quotient_32 <= _zz_rsp_payload_quotient_61[15:0];
    end else begin
      _zz_rsp_payload_quotient_32 <= _zz_rsp_payload_quotient_46[15:0];
    end
    _zz_rsp_payload_quotient_18 <= _zz_rsp_payload_quotient_17;
    _zz_rsp_payload_quotient_2 <= _zz__zz_rsp_payload_quotient_2[15:0];
    if(when_UnsignedDivider_l58_1) begin
      _zz_rsp_payload_quotient_33 <= _zz_rsp_payload_quotient_62[15:0];
    end else begin
      _zz_rsp_payload_quotient_33 <= _zz_rsp_payload_quotient_47[15:0];
    end
    _zz_rsp_payload_quotient_19 <= _zz_rsp_payload_quotient_18;
    _zz_rsp_payload_quotient_3 <= _zz__zz_rsp_payload_quotient_3[15:0];
    if(when_UnsignedDivider_l58_2) begin
      _zz_rsp_payload_quotient_34 <= _zz_rsp_payload_quotient_63[15:0];
    end else begin
      _zz_rsp_payload_quotient_34 <= _zz_rsp_payload_quotient_48[15:0];
    end
    _zz_rsp_payload_quotient_20 <= _zz_rsp_payload_quotient_19;
    _zz_rsp_payload_quotient_4 <= _zz__zz_rsp_payload_quotient_4[15:0];
    if(when_UnsignedDivider_l58_3) begin
      _zz_rsp_payload_quotient_35 <= _zz_rsp_payload_quotient_64[15:0];
    end else begin
      _zz_rsp_payload_quotient_35 <= _zz_rsp_payload_quotient_49[15:0];
    end
    _zz_rsp_payload_quotient_21 <= _zz_rsp_payload_quotient_20;
    _zz_rsp_payload_quotient_5 <= _zz__zz_rsp_payload_quotient_5[15:0];
    if(when_UnsignedDivider_l58_4) begin
      _zz_rsp_payload_quotient_36 <= _zz_rsp_payload_quotient_65[15:0];
    end else begin
      _zz_rsp_payload_quotient_36 <= _zz_rsp_payload_quotient_50[15:0];
    end
    _zz_rsp_payload_quotient_22 <= _zz_rsp_payload_quotient_21;
    _zz_rsp_payload_quotient_6 <= _zz__zz_rsp_payload_quotient_6[15:0];
    if(when_UnsignedDivider_l58_5) begin
      _zz_rsp_payload_quotient_37 <= _zz_rsp_payload_quotient_66[15:0];
    end else begin
      _zz_rsp_payload_quotient_37 <= _zz_rsp_payload_quotient_51[15:0];
    end
    _zz_rsp_payload_quotient_23 <= _zz_rsp_payload_quotient_22;
    _zz_rsp_payload_quotient_7 <= _zz__zz_rsp_payload_quotient_7[15:0];
    if(when_UnsignedDivider_l58_6) begin
      _zz_rsp_payload_quotient_38 <= _zz_rsp_payload_quotient_67[15:0];
    end else begin
      _zz_rsp_payload_quotient_38 <= _zz_rsp_payload_quotient_52[15:0];
    end
    _zz_rsp_payload_quotient_24 <= _zz_rsp_payload_quotient_23;
    _zz_rsp_payload_quotient_8 <= _zz__zz_rsp_payload_quotient_8[15:0];
    if(when_UnsignedDivider_l58_7) begin
      _zz_rsp_payload_quotient_39 <= _zz_rsp_payload_quotient_68[15:0];
    end else begin
      _zz_rsp_payload_quotient_39 <= _zz_rsp_payload_quotient_53[15:0];
    end
    _zz_rsp_payload_quotient_25 <= _zz_rsp_payload_quotient_24;
    _zz_rsp_payload_quotient_9 <= _zz__zz_rsp_payload_quotient_9[15:0];
    if(when_UnsignedDivider_l58_8) begin
      _zz_rsp_payload_quotient_40 <= _zz_rsp_payload_quotient_69[15:0];
    end else begin
      _zz_rsp_payload_quotient_40 <= _zz_rsp_payload_quotient_54[15:0];
    end
    _zz_rsp_payload_quotient_26 <= _zz_rsp_payload_quotient_25;
    _zz_rsp_payload_quotient_10 <= _zz__zz_rsp_payload_quotient_10[15:0];
    if(when_UnsignedDivider_l58_9) begin
      _zz_rsp_payload_quotient_41 <= _zz_rsp_payload_quotient_70[15:0];
    end else begin
      _zz_rsp_payload_quotient_41 <= _zz_rsp_payload_quotient_55[15:0];
    end
    _zz_rsp_payload_quotient_27 <= _zz_rsp_payload_quotient_26;
    _zz_rsp_payload_quotient_11 <= _zz__zz_rsp_payload_quotient_11[15:0];
    if(when_UnsignedDivider_l58_10) begin
      _zz_rsp_payload_quotient_42 <= _zz_rsp_payload_quotient_71[15:0];
    end else begin
      _zz_rsp_payload_quotient_42 <= _zz_rsp_payload_quotient_56[15:0];
    end
    _zz_rsp_payload_quotient_28 <= _zz_rsp_payload_quotient_27;
    _zz_rsp_payload_quotient_12 <= _zz__zz_rsp_payload_quotient_12[15:0];
    if(when_UnsignedDivider_l58_11) begin
      _zz_rsp_payload_quotient_43 <= _zz_rsp_payload_quotient_72[15:0];
    end else begin
      _zz_rsp_payload_quotient_43 <= _zz_rsp_payload_quotient_57[15:0];
    end
    _zz_rsp_payload_quotient_29 <= _zz_rsp_payload_quotient_28;
    _zz_rsp_payload_quotient_13 <= _zz__zz_rsp_payload_quotient_13[15:0];
    if(when_UnsignedDivider_l58_12) begin
      _zz_rsp_payload_quotient_44 <= _zz_rsp_payload_quotient_73[15:0];
    end else begin
      _zz_rsp_payload_quotient_44 <= _zz_rsp_payload_quotient_58[15:0];
    end
    _zz_rsp_payload_quotient_30 <= _zz_rsp_payload_quotient_29;
    _zz_rsp_payload_quotient_14 <= _zz__zz_rsp_payload_quotient_14[15:0];
    if(when_UnsignedDivider_l58_13) begin
      _zz_rsp_payload_quotient_45 <= _zz_rsp_payload_quotient_74[15:0];
    end else begin
      _zz_rsp_payload_quotient_45 <= _zz_rsp_payload_quotient_59[15:0];
    end
    _zz_rsp_payload_error <= _zz_rsp_payload_quotient_30;
    _zz_rsp_payload_quotient_15 <= _zz__zz_rsp_payload_quotient_15[15:0];
    if(when_UnsignedDivider_l58_14) begin
      _zz_rsp_payload_remainder <= _zz_rsp_payload_quotient_75[15:0];
    end else begin
      _zz_rsp_payload_remainder <= _zz_rsp_payload_quotient_60[15:0];
    end
  end


endmodule
