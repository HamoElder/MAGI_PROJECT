// Generator : SpinalHDL v1.6.0    git head : 73c8d8e2b86b45646e9d0b2e729291f2b65e6be3
// Component : OAMUnspinor
// Git hash  : 3aba5ba41129fa76a4728cd47203bcf10e3093cc



module OAMUnspinor (
  input               mod_iq_valid,
  output              mod_iq_ready,
  input      [15:0]   mod_iq_payload_cha_i,
  input      [15:0]   mod_iq_payload_cha_q,
  output              base_sub_iqs_valid,
  output     [31:0]   base_sub_iqs_payload_0_cha_i,
  output     [31:0]   base_sub_iqs_payload_0_cha_q,
  output     [31:0]   base_sub_iqs_payload_1_cha_i,
  output     [31:0]   base_sub_iqs_payload_1_cha_q,
  output     [31:0]   base_sub_iqs_payload_2_cha_i,
  output     [31:0]   base_sub_iqs_payload_2_cha_q,
  output     [31:0]   base_sub_iqs_payload_3_cha_i,
  output     [31:0]   base_sub_iqs_payload_3_cha_q,
  output     [31:0]   base_sub_iqs_payload_4_cha_i,
  output     [31:0]   base_sub_iqs_payload_4_cha_q,
  input               w_sel,
  input               w_en,
  input      [5:0]    w_addr,
  input      [15:0]   w_data,
  input               clk,
  input               resetn
);
  wire       [15:0]   oAMUnspin_5_shift_i_0;
  wire       [15:0]   oAMUnspin_5_shift_i_1;
  wire       [15:0]   oAMUnspin_5_shift_i_2;
  wire       [15:0]   oAMUnspin_5_shift_i_3;
  wire       [15:0]   oAMUnspin_5_shift_i_4;
  wire       [15:0]   oAMUnspin_5_shift_i_5;
  wire       [15:0]   oAMUnspin_5_shift_i_6;
  wire       [15:0]   oAMUnspin_5_shift_i_7;
  wire       [15:0]   oAMUnspin_5_shift_q_0;
  wire       [15:0]   oAMUnspin_5_shift_q_1;
  wire       [15:0]   oAMUnspin_5_shift_q_2;
  wire       [15:0]   oAMUnspin_5_shift_q_3;
  wire       [15:0]   oAMUnspin_5_shift_q_4;
  wire       [15:0]   oAMUnspin_5_shift_q_5;
  wire       [15:0]   oAMUnspin_5_shift_q_6;
  wire       [15:0]   oAMUnspin_5_shift_q_7;
  wire       [15:0]   oAMUnspin_6_shift_i_0;
  wire       [15:0]   oAMUnspin_6_shift_i_1;
  wire       [15:0]   oAMUnspin_6_shift_i_2;
  wire       [15:0]   oAMUnspin_6_shift_i_3;
  wire       [15:0]   oAMUnspin_6_shift_i_4;
  wire       [15:0]   oAMUnspin_6_shift_i_5;
  wire       [15:0]   oAMUnspin_6_shift_i_6;
  wire       [15:0]   oAMUnspin_6_shift_i_7;
  wire       [15:0]   oAMUnspin_6_shift_q_0;
  wire       [15:0]   oAMUnspin_6_shift_q_1;
  wire       [15:0]   oAMUnspin_6_shift_q_2;
  wire       [15:0]   oAMUnspin_6_shift_q_3;
  wire       [15:0]   oAMUnspin_6_shift_q_4;
  wire       [15:0]   oAMUnspin_6_shift_q_5;
  wire       [15:0]   oAMUnspin_6_shift_q_6;
  wire       [15:0]   oAMUnspin_6_shift_q_7;
  wire       [15:0]   oAMUnspin_7_shift_i_0;
  wire       [15:0]   oAMUnspin_7_shift_i_1;
  wire       [15:0]   oAMUnspin_7_shift_i_2;
  wire       [15:0]   oAMUnspin_7_shift_i_3;
  wire       [15:0]   oAMUnspin_7_shift_i_4;
  wire       [15:0]   oAMUnspin_7_shift_i_5;
  wire       [15:0]   oAMUnspin_7_shift_i_6;
  wire       [15:0]   oAMUnspin_7_shift_i_7;
  wire       [15:0]   oAMUnspin_7_shift_q_0;
  wire       [15:0]   oAMUnspin_7_shift_q_1;
  wire       [15:0]   oAMUnspin_7_shift_q_2;
  wire       [15:0]   oAMUnspin_7_shift_q_3;
  wire       [15:0]   oAMUnspin_7_shift_q_4;
  wire       [15:0]   oAMUnspin_7_shift_q_5;
  wire       [15:0]   oAMUnspin_7_shift_q_6;
  wire       [15:0]   oAMUnspin_7_shift_q_7;
  wire       [15:0]   oAMUnspin_8_shift_i_0;
  wire       [15:0]   oAMUnspin_8_shift_i_1;
  wire       [15:0]   oAMUnspin_8_shift_i_2;
  wire       [15:0]   oAMUnspin_8_shift_i_3;
  wire       [15:0]   oAMUnspin_8_shift_i_4;
  wire       [15:0]   oAMUnspin_8_shift_i_5;
  wire       [15:0]   oAMUnspin_8_shift_i_6;
  wire       [15:0]   oAMUnspin_8_shift_i_7;
  wire       [15:0]   oAMUnspin_8_shift_q_0;
  wire       [15:0]   oAMUnspin_8_shift_q_1;
  wire       [15:0]   oAMUnspin_8_shift_q_2;
  wire       [15:0]   oAMUnspin_8_shift_q_3;
  wire       [15:0]   oAMUnspin_8_shift_q_4;
  wire       [15:0]   oAMUnspin_8_shift_q_5;
  wire       [15:0]   oAMUnspin_8_shift_q_6;
  wire       [15:0]   oAMUnspin_8_shift_q_7;
  wire       [15:0]   oAMUnspin_9_shift_i_0;
  wire       [15:0]   oAMUnspin_9_shift_i_1;
  wire       [15:0]   oAMUnspin_9_shift_i_2;
  wire       [15:0]   oAMUnspin_9_shift_i_3;
  wire       [15:0]   oAMUnspin_9_shift_i_4;
  wire       [15:0]   oAMUnspin_9_shift_i_5;
  wire       [15:0]   oAMUnspin_9_shift_i_6;
  wire       [15:0]   oAMUnspin_9_shift_i_7;
  wire       [15:0]   oAMUnspin_9_shift_q_0;
  wire       [15:0]   oAMUnspin_9_shift_q_1;
  wire       [15:0]   oAMUnspin_9_shift_q_2;
  wire       [15:0]   oAMUnspin_9_shift_q_3;
  wire       [15:0]   oAMUnspin_9_shift_q_4;
  wire       [15:0]   oAMUnspin_9_shift_q_5;
  wire       [15:0]   oAMUnspin_9_shift_q_6;
  wire       [15:0]   oAMUnspin_9_shift_q_7;
  wire                oAMUnspin_5_base_sub_iq_valid;
  wire       [31:0]   oAMUnspin_5_base_sub_iq_payload_cha_i;
  wire       [31:0]   oAMUnspin_5_base_sub_iq_payload_cha_q;
  wire                oAMUnspin_6_base_sub_iq_valid;
  wire       [31:0]   oAMUnspin_6_base_sub_iq_payload_cha_i;
  wire       [31:0]   oAMUnspin_6_base_sub_iq_payload_cha_q;
  wire                oAMUnspin_7_base_sub_iq_valid;
  wire       [31:0]   oAMUnspin_7_base_sub_iq_payload_cha_i;
  wire       [31:0]   oAMUnspin_7_base_sub_iq_payload_cha_q;
  wire                oAMUnspin_8_base_sub_iq_valid;
  wire       [31:0]   oAMUnspin_8_base_sub_iq_payload_cha_i;
  wire       [31:0]   oAMUnspin_8_base_sub_iq_payload_cha_q;
  wire                oAMUnspin_9_base_sub_iq_valid;
  wire       [31:0]   oAMUnspin_9_base_sub_iq_payload_cha_i;
  wire       [31:0]   oAMUnspin_9_base_sub_iq_payload_cha_q;
  reg        [15:0]   _zz_shift_i_0;
  wire       [5:0]    _zz_shift_i_0_1;
  reg        [15:0]   _zz_shift_q_0;
  wire       [5:0]    _zz_shift_q_0_1;
  reg        [15:0]   _zz_shift_i_1;
  wire       [5:0]    _zz_shift_i_1_1;
  reg        [15:0]   _zz_shift_q_1;
  wire       [5:0]    _zz_shift_q_1_1;
  reg        [15:0]   _zz_shift_i_2;
  wire       [5:0]    _zz_shift_i_2_1;
  reg        [15:0]   _zz_shift_q_2;
  wire       [5:0]    _zz_shift_q_2_1;
  reg        [15:0]   _zz_shift_i_3;
  wire       [5:0]    _zz_shift_i_3_1;
  reg        [15:0]   _zz_shift_q_3;
  wire       [5:0]    _zz_shift_q_3_1;
  reg        [15:0]   _zz_shift_i_4;
  wire       [5:0]    _zz_shift_i_4_1;
  reg        [15:0]   _zz_shift_q_4;
  wire       [5:0]    _zz_shift_q_4_1;
  reg        [15:0]   _zz_shift_i_5;
  wire       [5:0]    _zz_shift_i_5_1;
  reg        [15:0]   _zz_shift_q_5;
  wire       [5:0]    _zz_shift_q_5_1;
  reg        [15:0]   _zz_shift_i_6;
  wire       [5:0]    _zz_shift_i_6_1;
  reg        [15:0]   _zz_shift_q_6;
  wire       [5:0]    _zz_shift_q_6_1;
  reg        [15:0]   _zz_shift_i_7;
  wire       [5:0]    _zz_shift_i_7_1;
  reg        [15:0]   _zz_shift_q_7;
  wire       [5:0]    _zz_shift_q_7_1;
  reg        [15:0]   _zz_shift_i_0_2;
  wire       [5:0]    _zz_shift_i_0_3;
  reg        [15:0]   _zz_shift_q_0_2;
  wire       [5:0]    _zz_shift_q_0_3;
  reg        [15:0]   _zz_shift_i_1_2;
  wire       [5:0]    _zz_shift_i_1_3;
  reg        [15:0]   _zz_shift_q_1_2;
  wire       [5:0]    _zz_shift_q_1_3;
  reg        [15:0]   _zz_shift_i_2_2;
  wire       [5:0]    _zz_shift_i_2_3;
  reg        [15:0]   _zz_shift_q_2_2;
  wire       [5:0]    _zz_shift_q_2_3;
  reg        [15:0]   _zz_shift_i_3_2;
  wire       [5:0]    _zz_shift_i_3_3;
  reg        [15:0]   _zz_shift_q_3_2;
  wire       [5:0]    _zz_shift_q_3_3;
  reg        [15:0]   _zz_shift_i_4_2;
  wire       [5:0]    _zz_shift_i_4_3;
  reg        [15:0]   _zz_shift_q_4_2;
  wire       [5:0]    _zz_shift_q_4_3;
  reg        [15:0]   _zz_shift_i_5_2;
  wire       [5:0]    _zz_shift_i_5_3;
  reg        [15:0]   _zz_shift_q_5_2;
  wire       [5:0]    _zz_shift_q_5_3;
  reg        [15:0]   _zz_shift_i_6_2;
  wire       [5:0]    _zz_shift_i_6_3;
  reg        [15:0]   _zz_shift_q_6_2;
  wire       [5:0]    _zz_shift_q_6_3;
  reg        [15:0]   _zz_shift_i_7_2;
  wire       [5:0]    _zz_shift_i_7_3;
  reg        [15:0]   _zz_shift_q_7_2;
  wire       [5:0]    _zz_shift_q_7_3;
  reg        [15:0]   _zz_shift_i_0_4;
  wire       [5:0]    _zz_shift_i_0_5;
  reg        [15:0]   _zz_shift_q_0_4;
  wire       [5:0]    _zz_shift_q_0_5;
  reg        [15:0]   _zz_shift_i_1_4;
  wire       [5:0]    _zz_shift_i_1_5;
  reg        [15:0]   _zz_shift_q_1_4;
  wire       [5:0]    _zz_shift_q_1_5;
  reg        [15:0]   _zz_shift_i_2_4;
  wire       [5:0]    _zz_shift_i_2_5;
  reg        [15:0]   _zz_shift_q_2_4;
  wire       [5:0]    _zz_shift_q_2_5;
  reg        [15:0]   _zz_shift_i_3_4;
  wire       [5:0]    _zz_shift_i_3_5;
  reg        [15:0]   _zz_shift_q_3_4;
  wire       [5:0]    _zz_shift_q_3_5;
  reg        [15:0]   _zz_shift_i_4_4;
  wire       [5:0]    _zz_shift_i_4_5;
  reg        [15:0]   _zz_shift_q_4_4;
  wire       [5:0]    _zz_shift_q_4_5;
  reg        [15:0]   _zz_shift_i_5_4;
  wire       [5:0]    _zz_shift_i_5_5;
  reg        [15:0]   _zz_shift_q_5_4;
  wire       [5:0]    _zz_shift_q_5_5;
  reg        [15:0]   _zz_shift_i_6_4;
  wire       [5:0]    _zz_shift_i_6_5;
  reg        [15:0]   _zz_shift_q_6_4;
  wire       [5:0]    _zz_shift_q_6_5;
  reg        [15:0]   _zz_shift_i_7_4;
  wire       [5:0]    _zz_shift_i_7_5;
  reg        [15:0]   _zz_shift_q_7_4;
  wire       [5:0]    _zz_shift_q_7_5;
  reg        [15:0]   _zz_shift_i_0_6;
  wire       [5:0]    _zz_shift_i_0_7;
  reg        [15:0]   _zz_shift_q_0_6;
  wire       [5:0]    _zz_shift_q_0_7;
  reg        [15:0]   _zz_shift_i_1_6;
  wire       [5:0]    _zz_shift_i_1_7;
  reg        [15:0]   _zz_shift_q_1_6;
  wire       [5:0]    _zz_shift_q_1_7;
  reg        [15:0]   _zz_shift_i_2_6;
  wire       [5:0]    _zz_shift_i_2_7;
  reg        [15:0]   _zz_shift_q_2_6;
  wire       [5:0]    _zz_shift_q_2_7;
  reg        [15:0]   _zz_shift_i_3_6;
  wire       [5:0]    _zz_shift_i_3_7;
  reg        [15:0]   _zz_shift_q_3_6;
  wire       [5:0]    _zz_shift_q_3_7;
  reg        [15:0]   _zz_shift_i_4_6;
  wire       [5:0]    _zz_shift_i_4_7;
  reg        [15:0]   _zz_shift_q_4_6;
  wire       [5:0]    _zz_shift_q_4_7;
  reg        [15:0]   _zz_shift_i_5_6;
  wire       [5:0]    _zz_shift_i_5_7;
  reg        [15:0]   _zz_shift_q_5_6;
  wire       [5:0]    _zz_shift_q_5_7;
  reg        [15:0]   _zz_shift_i_6_6;
  wire       [5:0]    _zz_shift_i_6_7;
  reg        [15:0]   _zz_shift_q_6_6;
  wire       [5:0]    _zz_shift_q_6_7;
  reg        [15:0]   _zz_shift_i_7_6;
  wire       [5:0]    _zz_shift_i_7_7;
  reg        [15:0]   _zz_shift_q_7_6;
  wire       [5:0]    _zz_shift_q_7_7;
  reg        [15:0]   _zz_shift_i_0_8;
  wire       [5:0]    _zz_shift_i_0_9;
  reg        [15:0]   _zz_shift_q_0_8;
  wire       [5:0]    _zz_shift_q_0_9;
  reg        [15:0]   _zz_shift_i_1_8;
  wire       [5:0]    _zz_shift_i_1_9;
  reg        [15:0]   _zz_shift_q_1_8;
  wire       [5:0]    _zz_shift_q_1_9;
  reg        [15:0]   _zz_shift_i_2_8;
  wire       [5:0]    _zz_shift_i_2_9;
  reg        [15:0]   _zz_shift_q_2_8;
  wire       [5:0]    _zz_shift_q_2_9;
  reg        [15:0]   _zz_shift_i_3_8;
  wire       [5:0]    _zz_shift_i_3_9;
  reg        [15:0]   _zz_shift_q_3_8;
  wire       [5:0]    _zz_shift_q_3_9;
  reg        [15:0]   _zz_shift_i_4_8;
  wire       [5:0]    _zz_shift_i_4_9;
  reg        [15:0]   _zz_shift_q_4_8;
  wire       [5:0]    _zz_shift_q_4_9;
  reg        [15:0]   _zz_shift_i_5_8;
  wire       [5:0]    _zz_shift_i_5_9;
  reg        [15:0]   _zz_shift_q_5_8;
  wire       [5:0]    _zz_shift_q_5_9;
  reg        [15:0]   _zz_shift_i_6_8;
  wire       [5:0]    _zz_shift_i_6_9;
  reg        [15:0]   _zz_shift_q_6_8;
  wire       [5:0]    _zz_shift_q_6_9;
  reg        [15:0]   _zz_shift_i_7_8;
  wire       [5:0]    _zz_shift_i_7_9;
  reg        [15:0]   _zz_shift_q_7_8;
  wire       [5:0]    _zz_shift_q_7_9;
  reg        [15:0]   shift_i_map_0;
  reg        [15:0]   shift_i_map_1;
  reg        [15:0]   shift_i_map_2;
  reg        [15:0]   shift_i_map_3;
  reg        [15:0]   shift_i_map_4;
  reg        [15:0]   shift_i_map_5;
  reg        [15:0]   shift_i_map_6;
  reg        [15:0]   shift_i_map_7;
  reg        [15:0]   shift_i_map_8;
  reg        [15:0]   shift_i_map_9;
  reg        [15:0]   shift_i_map_10;
  reg        [15:0]   shift_i_map_11;
  reg        [15:0]   shift_i_map_12;
  reg        [15:0]   shift_i_map_13;
  reg        [15:0]   shift_i_map_14;
  reg        [15:0]   shift_i_map_15;
  reg        [15:0]   shift_i_map_16;
  reg        [15:0]   shift_i_map_17;
  reg        [15:0]   shift_i_map_18;
  reg        [15:0]   shift_i_map_19;
  reg        [15:0]   shift_i_map_20;
  reg        [15:0]   shift_i_map_21;
  reg        [15:0]   shift_i_map_22;
  reg        [15:0]   shift_i_map_23;
  reg        [15:0]   shift_i_map_24;
  reg        [15:0]   shift_i_map_25;
  reg        [15:0]   shift_i_map_26;
  reg        [15:0]   shift_i_map_27;
  reg        [15:0]   shift_i_map_28;
  reg        [15:0]   shift_i_map_29;
  reg        [15:0]   shift_i_map_30;
  reg        [15:0]   shift_i_map_31;
  reg        [15:0]   shift_i_map_32;
  reg        [15:0]   shift_i_map_33;
  reg        [15:0]   shift_i_map_34;
  reg        [15:0]   shift_i_map_35;
  reg        [15:0]   shift_i_map_36;
  reg        [15:0]   shift_i_map_37;
  reg        [15:0]   shift_i_map_38;
  reg        [15:0]   shift_i_map_39;
  reg        [15:0]   shift_q_map_0;
  reg        [15:0]   shift_q_map_1;
  reg        [15:0]   shift_q_map_2;
  reg        [15:0]   shift_q_map_3;
  reg        [15:0]   shift_q_map_4;
  reg        [15:0]   shift_q_map_5;
  reg        [15:0]   shift_q_map_6;
  reg        [15:0]   shift_q_map_7;
  reg        [15:0]   shift_q_map_8;
  reg        [15:0]   shift_q_map_9;
  reg        [15:0]   shift_q_map_10;
  reg        [15:0]   shift_q_map_11;
  reg        [15:0]   shift_q_map_12;
  reg        [15:0]   shift_q_map_13;
  reg        [15:0]   shift_q_map_14;
  reg        [15:0]   shift_q_map_15;
  reg        [15:0]   shift_q_map_16;
  reg        [15:0]   shift_q_map_17;
  reg        [15:0]   shift_q_map_18;
  reg        [15:0]   shift_q_map_19;
  reg        [15:0]   shift_q_map_20;
  reg        [15:0]   shift_q_map_21;
  reg        [15:0]   shift_q_map_22;
  reg        [15:0]   shift_q_map_23;
  reg        [15:0]   shift_q_map_24;
  reg        [15:0]   shift_q_map_25;
  reg        [15:0]   shift_q_map_26;
  reg        [15:0]   shift_q_map_27;
  reg        [15:0]   shift_q_map_28;
  reg        [15:0]   shift_q_map_29;
  reg        [15:0]   shift_q_map_30;
  reg        [15:0]   shift_q_map_31;
  reg        [15:0]   shift_q_map_32;
  reg        [15:0]   shift_q_map_33;
  reg        [15:0]   shift_q_map_34;
  reg        [15:0]   shift_q_map_35;
  reg        [15:0]   shift_q_map_36;
  reg        [15:0]   shift_q_map_37;
  reg        [15:0]   shift_q_map_38;
  reg        [15:0]   shift_q_map_39;
  wire       [63:0]   _zz_1;
  wire       [63:0]   _zz_2;
  wire                base_sub_valid_vec_0;
  wire                base_sub_valid_vec_1;
  wire                base_sub_valid_vec_2;
  wire                base_sub_valid_vec_3;
  wire                base_sub_valid_vec_4;

  assign _zz_shift_i_0_1 = 6'h0;
  assign _zz_shift_q_0_1 = 6'h0;
  assign _zz_shift_i_1_1 = 6'h01;
  assign _zz_shift_q_1_1 = 6'h01;
  assign _zz_shift_i_2_1 = 6'h02;
  assign _zz_shift_q_2_1 = 6'h02;
  assign _zz_shift_i_3_1 = 6'h03;
  assign _zz_shift_q_3_1 = 6'h03;
  assign _zz_shift_i_4_1 = 6'h04;
  assign _zz_shift_q_4_1 = 6'h04;
  assign _zz_shift_i_5_1 = 6'h05;
  assign _zz_shift_q_5_1 = 6'h05;
  assign _zz_shift_i_6_1 = 6'h06;
  assign _zz_shift_q_6_1 = 6'h06;
  assign _zz_shift_i_7_1 = 6'h07;
  assign _zz_shift_q_7_1 = 6'h07;
  assign _zz_shift_i_0_3 = 6'h08;
  assign _zz_shift_q_0_3 = 6'h08;
  assign _zz_shift_i_1_3 = 6'h09;
  assign _zz_shift_q_1_3 = 6'h09;
  assign _zz_shift_i_2_3 = 6'h0a;
  assign _zz_shift_q_2_3 = 6'h0a;
  assign _zz_shift_i_3_3 = 6'h0b;
  assign _zz_shift_q_3_3 = 6'h0b;
  assign _zz_shift_i_4_3 = 6'h0c;
  assign _zz_shift_q_4_3 = 6'h0c;
  assign _zz_shift_i_5_3 = 6'h0d;
  assign _zz_shift_q_5_3 = 6'h0d;
  assign _zz_shift_i_6_3 = 6'h0e;
  assign _zz_shift_q_6_3 = 6'h0e;
  assign _zz_shift_i_7_3 = 6'h0f;
  assign _zz_shift_q_7_3 = 6'h0f;
  assign _zz_shift_i_0_5 = 6'h10;
  assign _zz_shift_q_0_5 = 6'h10;
  assign _zz_shift_i_1_5 = 6'h11;
  assign _zz_shift_q_1_5 = 6'h11;
  assign _zz_shift_i_2_5 = 6'h12;
  assign _zz_shift_q_2_5 = 6'h12;
  assign _zz_shift_i_3_5 = 6'h13;
  assign _zz_shift_q_3_5 = 6'h13;
  assign _zz_shift_i_4_5 = 6'h14;
  assign _zz_shift_q_4_5 = 6'h14;
  assign _zz_shift_i_5_5 = 6'h15;
  assign _zz_shift_q_5_5 = 6'h15;
  assign _zz_shift_i_6_5 = 6'h16;
  assign _zz_shift_q_6_5 = 6'h16;
  assign _zz_shift_i_7_5 = 6'h17;
  assign _zz_shift_q_7_5 = 6'h17;
  assign _zz_shift_i_0_7 = 6'h18;
  assign _zz_shift_q_0_7 = 6'h18;
  assign _zz_shift_i_1_7 = 6'h19;
  assign _zz_shift_q_1_7 = 6'h19;
  assign _zz_shift_i_2_7 = 6'h1a;
  assign _zz_shift_q_2_7 = 6'h1a;
  assign _zz_shift_i_3_7 = 6'h1b;
  assign _zz_shift_q_3_7 = 6'h1b;
  assign _zz_shift_i_4_7 = 6'h1c;
  assign _zz_shift_q_4_7 = 6'h1c;
  assign _zz_shift_i_5_7 = 6'h1d;
  assign _zz_shift_q_5_7 = 6'h1d;
  assign _zz_shift_i_6_7 = 6'h1e;
  assign _zz_shift_q_6_7 = 6'h1e;
  assign _zz_shift_i_7_7 = 6'h1f;
  assign _zz_shift_q_7_7 = 6'h1f;
  assign _zz_shift_i_0_9 = 6'h20;
  assign _zz_shift_q_0_9 = 6'h20;
  assign _zz_shift_i_1_9 = 6'h21;
  assign _zz_shift_q_1_9 = 6'h21;
  assign _zz_shift_i_2_9 = 6'h22;
  assign _zz_shift_q_2_9 = 6'h22;
  assign _zz_shift_i_3_9 = 6'h23;
  assign _zz_shift_q_3_9 = 6'h23;
  assign _zz_shift_i_4_9 = 6'h24;
  assign _zz_shift_q_4_9 = 6'h24;
  assign _zz_shift_i_5_9 = 6'h25;
  assign _zz_shift_q_5_9 = 6'h25;
  assign _zz_shift_i_6_9 = 6'h26;
  assign _zz_shift_q_6_9 = 6'h26;
  assign _zz_shift_i_7_9 = 6'h27;
  assign _zz_shift_q_7_9 = 6'h27;
  OAMUnspin oAMUnspin_5 (
    .shift_i_0                    (oAMUnspin_5_shift_i_0                  ), //i
    .shift_i_1                    (oAMUnspin_5_shift_i_1                  ), //i
    .shift_i_2                    (oAMUnspin_5_shift_i_2                  ), //i
    .shift_i_3                    (oAMUnspin_5_shift_i_3                  ), //i
    .shift_i_4                    (oAMUnspin_5_shift_i_4                  ), //i
    .shift_i_5                    (oAMUnspin_5_shift_i_5                  ), //i
    .shift_i_6                    (oAMUnspin_5_shift_i_6                  ), //i
    .shift_i_7                    (oAMUnspin_5_shift_i_7                  ), //i
    .shift_q_0                    (oAMUnspin_5_shift_q_0                  ), //i
    .shift_q_1                    (oAMUnspin_5_shift_q_1                  ), //i
    .shift_q_2                    (oAMUnspin_5_shift_q_2                  ), //i
    .shift_q_3                    (oAMUnspin_5_shift_q_3                  ), //i
    .shift_q_4                    (oAMUnspin_5_shift_q_4                  ), //i
    .shift_q_5                    (oAMUnspin_5_shift_q_5                  ), //i
    .shift_q_6                    (oAMUnspin_5_shift_q_6                  ), //i
    .shift_q_7                    (oAMUnspin_5_shift_q_7                  ), //i
    .mod_iq_valid                 (mod_iq_valid                           ), //i
    .mod_iq_payload_cha_i         (mod_iq_payload_cha_i                   ), //i
    .mod_iq_payload_cha_q         (mod_iq_payload_cha_q                   ), //i
    .base_sub_iq_valid            (oAMUnspin_5_base_sub_iq_valid          ), //o
    .base_sub_iq_payload_cha_i    (oAMUnspin_5_base_sub_iq_payload_cha_i  ), //o
    .base_sub_iq_payload_cha_q    (oAMUnspin_5_base_sub_iq_payload_cha_q  ), //o
    .clk                          (clk                                    ), //i
    .resetn                       (resetn                                 )  //i
  );
  OAMUnspin oAMUnspin_6 (
    .shift_i_0                    (oAMUnspin_6_shift_i_0                  ), //i
    .shift_i_1                    (oAMUnspin_6_shift_i_1                  ), //i
    .shift_i_2                    (oAMUnspin_6_shift_i_2                  ), //i
    .shift_i_3                    (oAMUnspin_6_shift_i_3                  ), //i
    .shift_i_4                    (oAMUnspin_6_shift_i_4                  ), //i
    .shift_i_5                    (oAMUnspin_6_shift_i_5                  ), //i
    .shift_i_6                    (oAMUnspin_6_shift_i_6                  ), //i
    .shift_i_7                    (oAMUnspin_6_shift_i_7                  ), //i
    .shift_q_0                    (oAMUnspin_6_shift_q_0                  ), //i
    .shift_q_1                    (oAMUnspin_6_shift_q_1                  ), //i
    .shift_q_2                    (oAMUnspin_6_shift_q_2                  ), //i
    .shift_q_3                    (oAMUnspin_6_shift_q_3                  ), //i
    .shift_q_4                    (oAMUnspin_6_shift_q_4                  ), //i
    .shift_q_5                    (oAMUnspin_6_shift_q_5                  ), //i
    .shift_q_6                    (oAMUnspin_6_shift_q_6                  ), //i
    .shift_q_7                    (oAMUnspin_6_shift_q_7                  ), //i
    .mod_iq_valid                 (mod_iq_valid                           ), //i
    .mod_iq_payload_cha_i         (mod_iq_payload_cha_i                   ), //i
    .mod_iq_payload_cha_q         (mod_iq_payload_cha_q                   ), //i
    .base_sub_iq_valid            (oAMUnspin_6_base_sub_iq_valid          ), //o
    .base_sub_iq_payload_cha_i    (oAMUnspin_6_base_sub_iq_payload_cha_i  ), //o
    .base_sub_iq_payload_cha_q    (oAMUnspin_6_base_sub_iq_payload_cha_q  ), //o
    .clk                          (clk                                    ), //i
    .resetn                       (resetn                                 )  //i
  );
  OAMUnspin oAMUnspin_7 (
    .shift_i_0                    (oAMUnspin_7_shift_i_0                  ), //i
    .shift_i_1                    (oAMUnspin_7_shift_i_1                  ), //i
    .shift_i_2                    (oAMUnspin_7_shift_i_2                  ), //i
    .shift_i_3                    (oAMUnspin_7_shift_i_3                  ), //i
    .shift_i_4                    (oAMUnspin_7_shift_i_4                  ), //i
    .shift_i_5                    (oAMUnspin_7_shift_i_5                  ), //i
    .shift_i_6                    (oAMUnspin_7_shift_i_6                  ), //i
    .shift_i_7                    (oAMUnspin_7_shift_i_7                  ), //i
    .shift_q_0                    (oAMUnspin_7_shift_q_0                  ), //i
    .shift_q_1                    (oAMUnspin_7_shift_q_1                  ), //i
    .shift_q_2                    (oAMUnspin_7_shift_q_2                  ), //i
    .shift_q_3                    (oAMUnspin_7_shift_q_3                  ), //i
    .shift_q_4                    (oAMUnspin_7_shift_q_4                  ), //i
    .shift_q_5                    (oAMUnspin_7_shift_q_5                  ), //i
    .shift_q_6                    (oAMUnspin_7_shift_q_6                  ), //i
    .shift_q_7                    (oAMUnspin_7_shift_q_7                  ), //i
    .mod_iq_valid                 (mod_iq_valid                           ), //i
    .mod_iq_payload_cha_i         (mod_iq_payload_cha_i                   ), //i
    .mod_iq_payload_cha_q         (mod_iq_payload_cha_q                   ), //i
    .base_sub_iq_valid            (oAMUnspin_7_base_sub_iq_valid          ), //o
    .base_sub_iq_payload_cha_i    (oAMUnspin_7_base_sub_iq_payload_cha_i  ), //o
    .base_sub_iq_payload_cha_q    (oAMUnspin_7_base_sub_iq_payload_cha_q  ), //o
    .clk                          (clk                                    ), //i
    .resetn                       (resetn                                 )  //i
  );
  OAMUnspin oAMUnspin_8 (
    .shift_i_0                    (oAMUnspin_8_shift_i_0                  ), //i
    .shift_i_1                    (oAMUnspin_8_shift_i_1                  ), //i
    .shift_i_2                    (oAMUnspin_8_shift_i_2                  ), //i
    .shift_i_3                    (oAMUnspin_8_shift_i_3                  ), //i
    .shift_i_4                    (oAMUnspin_8_shift_i_4                  ), //i
    .shift_i_5                    (oAMUnspin_8_shift_i_5                  ), //i
    .shift_i_6                    (oAMUnspin_8_shift_i_6                  ), //i
    .shift_i_7                    (oAMUnspin_8_shift_i_7                  ), //i
    .shift_q_0                    (oAMUnspin_8_shift_q_0                  ), //i
    .shift_q_1                    (oAMUnspin_8_shift_q_1                  ), //i
    .shift_q_2                    (oAMUnspin_8_shift_q_2                  ), //i
    .shift_q_3                    (oAMUnspin_8_shift_q_3                  ), //i
    .shift_q_4                    (oAMUnspin_8_shift_q_4                  ), //i
    .shift_q_5                    (oAMUnspin_8_shift_q_5                  ), //i
    .shift_q_6                    (oAMUnspin_8_shift_q_6                  ), //i
    .shift_q_7                    (oAMUnspin_8_shift_q_7                  ), //i
    .mod_iq_valid                 (mod_iq_valid                           ), //i
    .mod_iq_payload_cha_i         (mod_iq_payload_cha_i                   ), //i
    .mod_iq_payload_cha_q         (mod_iq_payload_cha_q                   ), //i
    .base_sub_iq_valid            (oAMUnspin_8_base_sub_iq_valid          ), //o
    .base_sub_iq_payload_cha_i    (oAMUnspin_8_base_sub_iq_payload_cha_i  ), //o
    .base_sub_iq_payload_cha_q    (oAMUnspin_8_base_sub_iq_payload_cha_q  ), //o
    .clk                          (clk                                    ), //i
    .resetn                       (resetn                                 )  //i
  );
  OAMUnspin oAMUnspin_9 (
    .shift_i_0                    (oAMUnspin_9_shift_i_0                  ), //i
    .shift_i_1                    (oAMUnspin_9_shift_i_1                  ), //i
    .shift_i_2                    (oAMUnspin_9_shift_i_2                  ), //i
    .shift_i_3                    (oAMUnspin_9_shift_i_3                  ), //i
    .shift_i_4                    (oAMUnspin_9_shift_i_4                  ), //i
    .shift_i_5                    (oAMUnspin_9_shift_i_5                  ), //i
    .shift_i_6                    (oAMUnspin_9_shift_i_6                  ), //i
    .shift_i_7                    (oAMUnspin_9_shift_i_7                  ), //i
    .shift_q_0                    (oAMUnspin_9_shift_q_0                  ), //i
    .shift_q_1                    (oAMUnspin_9_shift_q_1                  ), //i
    .shift_q_2                    (oAMUnspin_9_shift_q_2                  ), //i
    .shift_q_3                    (oAMUnspin_9_shift_q_3                  ), //i
    .shift_q_4                    (oAMUnspin_9_shift_q_4                  ), //i
    .shift_q_5                    (oAMUnspin_9_shift_q_5                  ), //i
    .shift_q_6                    (oAMUnspin_9_shift_q_6                  ), //i
    .shift_q_7                    (oAMUnspin_9_shift_q_7                  ), //i
    .mod_iq_valid                 (mod_iq_valid                           ), //i
    .mod_iq_payload_cha_i         (mod_iq_payload_cha_i                   ), //i
    .mod_iq_payload_cha_q         (mod_iq_payload_cha_q                   ), //i
    .base_sub_iq_valid            (oAMUnspin_9_base_sub_iq_valid          ), //o
    .base_sub_iq_payload_cha_i    (oAMUnspin_9_base_sub_iq_payload_cha_i  ), //o
    .base_sub_iq_payload_cha_q    (oAMUnspin_9_base_sub_iq_payload_cha_q  ), //o
    .clk                          (clk                                    ), //i
    .resetn                       (resetn                                 )  //i
  );
  always @(*) begin
    case(_zz_shift_i_0_1)
      6'b000000 : begin
        _zz_shift_i_0 = shift_i_map_0;
      end
      6'b000001 : begin
        _zz_shift_i_0 = shift_i_map_1;
      end
      6'b000010 : begin
        _zz_shift_i_0 = shift_i_map_2;
      end
      6'b000011 : begin
        _zz_shift_i_0 = shift_i_map_3;
      end
      6'b000100 : begin
        _zz_shift_i_0 = shift_i_map_4;
      end
      6'b000101 : begin
        _zz_shift_i_0 = shift_i_map_5;
      end
      6'b000110 : begin
        _zz_shift_i_0 = shift_i_map_6;
      end
      6'b000111 : begin
        _zz_shift_i_0 = shift_i_map_7;
      end
      6'b001000 : begin
        _zz_shift_i_0 = shift_i_map_8;
      end
      6'b001001 : begin
        _zz_shift_i_0 = shift_i_map_9;
      end
      6'b001010 : begin
        _zz_shift_i_0 = shift_i_map_10;
      end
      6'b001011 : begin
        _zz_shift_i_0 = shift_i_map_11;
      end
      6'b001100 : begin
        _zz_shift_i_0 = shift_i_map_12;
      end
      6'b001101 : begin
        _zz_shift_i_0 = shift_i_map_13;
      end
      6'b001110 : begin
        _zz_shift_i_0 = shift_i_map_14;
      end
      6'b001111 : begin
        _zz_shift_i_0 = shift_i_map_15;
      end
      6'b010000 : begin
        _zz_shift_i_0 = shift_i_map_16;
      end
      6'b010001 : begin
        _zz_shift_i_0 = shift_i_map_17;
      end
      6'b010010 : begin
        _zz_shift_i_0 = shift_i_map_18;
      end
      6'b010011 : begin
        _zz_shift_i_0 = shift_i_map_19;
      end
      6'b010100 : begin
        _zz_shift_i_0 = shift_i_map_20;
      end
      6'b010101 : begin
        _zz_shift_i_0 = shift_i_map_21;
      end
      6'b010110 : begin
        _zz_shift_i_0 = shift_i_map_22;
      end
      6'b010111 : begin
        _zz_shift_i_0 = shift_i_map_23;
      end
      6'b011000 : begin
        _zz_shift_i_0 = shift_i_map_24;
      end
      6'b011001 : begin
        _zz_shift_i_0 = shift_i_map_25;
      end
      6'b011010 : begin
        _zz_shift_i_0 = shift_i_map_26;
      end
      6'b011011 : begin
        _zz_shift_i_0 = shift_i_map_27;
      end
      6'b011100 : begin
        _zz_shift_i_0 = shift_i_map_28;
      end
      6'b011101 : begin
        _zz_shift_i_0 = shift_i_map_29;
      end
      6'b011110 : begin
        _zz_shift_i_0 = shift_i_map_30;
      end
      6'b011111 : begin
        _zz_shift_i_0 = shift_i_map_31;
      end
      6'b100000 : begin
        _zz_shift_i_0 = shift_i_map_32;
      end
      6'b100001 : begin
        _zz_shift_i_0 = shift_i_map_33;
      end
      6'b100010 : begin
        _zz_shift_i_0 = shift_i_map_34;
      end
      6'b100011 : begin
        _zz_shift_i_0 = shift_i_map_35;
      end
      6'b100100 : begin
        _zz_shift_i_0 = shift_i_map_36;
      end
      6'b100101 : begin
        _zz_shift_i_0 = shift_i_map_37;
      end
      6'b100110 : begin
        _zz_shift_i_0 = shift_i_map_38;
      end
      default : begin
        _zz_shift_i_0 = shift_i_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_0_1)
      6'b000000 : begin
        _zz_shift_q_0 = shift_q_map_0;
      end
      6'b000001 : begin
        _zz_shift_q_0 = shift_q_map_1;
      end
      6'b000010 : begin
        _zz_shift_q_0 = shift_q_map_2;
      end
      6'b000011 : begin
        _zz_shift_q_0 = shift_q_map_3;
      end
      6'b000100 : begin
        _zz_shift_q_0 = shift_q_map_4;
      end
      6'b000101 : begin
        _zz_shift_q_0 = shift_q_map_5;
      end
      6'b000110 : begin
        _zz_shift_q_0 = shift_q_map_6;
      end
      6'b000111 : begin
        _zz_shift_q_0 = shift_q_map_7;
      end
      6'b001000 : begin
        _zz_shift_q_0 = shift_q_map_8;
      end
      6'b001001 : begin
        _zz_shift_q_0 = shift_q_map_9;
      end
      6'b001010 : begin
        _zz_shift_q_0 = shift_q_map_10;
      end
      6'b001011 : begin
        _zz_shift_q_0 = shift_q_map_11;
      end
      6'b001100 : begin
        _zz_shift_q_0 = shift_q_map_12;
      end
      6'b001101 : begin
        _zz_shift_q_0 = shift_q_map_13;
      end
      6'b001110 : begin
        _zz_shift_q_0 = shift_q_map_14;
      end
      6'b001111 : begin
        _zz_shift_q_0 = shift_q_map_15;
      end
      6'b010000 : begin
        _zz_shift_q_0 = shift_q_map_16;
      end
      6'b010001 : begin
        _zz_shift_q_0 = shift_q_map_17;
      end
      6'b010010 : begin
        _zz_shift_q_0 = shift_q_map_18;
      end
      6'b010011 : begin
        _zz_shift_q_0 = shift_q_map_19;
      end
      6'b010100 : begin
        _zz_shift_q_0 = shift_q_map_20;
      end
      6'b010101 : begin
        _zz_shift_q_0 = shift_q_map_21;
      end
      6'b010110 : begin
        _zz_shift_q_0 = shift_q_map_22;
      end
      6'b010111 : begin
        _zz_shift_q_0 = shift_q_map_23;
      end
      6'b011000 : begin
        _zz_shift_q_0 = shift_q_map_24;
      end
      6'b011001 : begin
        _zz_shift_q_0 = shift_q_map_25;
      end
      6'b011010 : begin
        _zz_shift_q_0 = shift_q_map_26;
      end
      6'b011011 : begin
        _zz_shift_q_0 = shift_q_map_27;
      end
      6'b011100 : begin
        _zz_shift_q_0 = shift_q_map_28;
      end
      6'b011101 : begin
        _zz_shift_q_0 = shift_q_map_29;
      end
      6'b011110 : begin
        _zz_shift_q_0 = shift_q_map_30;
      end
      6'b011111 : begin
        _zz_shift_q_0 = shift_q_map_31;
      end
      6'b100000 : begin
        _zz_shift_q_0 = shift_q_map_32;
      end
      6'b100001 : begin
        _zz_shift_q_0 = shift_q_map_33;
      end
      6'b100010 : begin
        _zz_shift_q_0 = shift_q_map_34;
      end
      6'b100011 : begin
        _zz_shift_q_0 = shift_q_map_35;
      end
      6'b100100 : begin
        _zz_shift_q_0 = shift_q_map_36;
      end
      6'b100101 : begin
        _zz_shift_q_0 = shift_q_map_37;
      end
      6'b100110 : begin
        _zz_shift_q_0 = shift_q_map_38;
      end
      default : begin
        _zz_shift_q_0 = shift_q_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_1_1)
      6'b000000 : begin
        _zz_shift_i_1 = shift_i_map_0;
      end
      6'b000001 : begin
        _zz_shift_i_1 = shift_i_map_1;
      end
      6'b000010 : begin
        _zz_shift_i_1 = shift_i_map_2;
      end
      6'b000011 : begin
        _zz_shift_i_1 = shift_i_map_3;
      end
      6'b000100 : begin
        _zz_shift_i_1 = shift_i_map_4;
      end
      6'b000101 : begin
        _zz_shift_i_1 = shift_i_map_5;
      end
      6'b000110 : begin
        _zz_shift_i_1 = shift_i_map_6;
      end
      6'b000111 : begin
        _zz_shift_i_1 = shift_i_map_7;
      end
      6'b001000 : begin
        _zz_shift_i_1 = shift_i_map_8;
      end
      6'b001001 : begin
        _zz_shift_i_1 = shift_i_map_9;
      end
      6'b001010 : begin
        _zz_shift_i_1 = shift_i_map_10;
      end
      6'b001011 : begin
        _zz_shift_i_1 = shift_i_map_11;
      end
      6'b001100 : begin
        _zz_shift_i_1 = shift_i_map_12;
      end
      6'b001101 : begin
        _zz_shift_i_1 = shift_i_map_13;
      end
      6'b001110 : begin
        _zz_shift_i_1 = shift_i_map_14;
      end
      6'b001111 : begin
        _zz_shift_i_1 = shift_i_map_15;
      end
      6'b010000 : begin
        _zz_shift_i_1 = shift_i_map_16;
      end
      6'b010001 : begin
        _zz_shift_i_1 = shift_i_map_17;
      end
      6'b010010 : begin
        _zz_shift_i_1 = shift_i_map_18;
      end
      6'b010011 : begin
        _zz_shift_i_1 = shift_i_map_19;
      end
      6'b010100 : begin
        _zz_shift_i_1 = shift_i_map_20;
      end
      6'b010101 : begin
        _zz_shift_i_1 = shift_i_map_21;
      end
      6'b010110 : begin
        _zz_shift_i_1 = shift_i_map_22;
      end
      6'b010111 : begin
        _zz_shift_i_1 = shift_i_map_23;
      end
      6'b011000 : begin
        _zz_shift_i_1 = shift_i_map_24;
      end
      6'b011001 : begin
        _zz_shift_i_1 = shift_i_map_25;
      end
      6'b011010 : begin
        _zz_shift_i_1 = shift_i_map_26;
      end
      6'b011011 : begin
        _zz_shift_i_1 = shift_i_map_27;
      end
      6'b011100 : begin
        _zz_shift_i_1 = shift_i_map_28;
      end
      6'b011101 : begin
        _zz_shift_i_1 = shift_i_map_29;
      end
      6'b011110 : begin
        _zz_shift_i_1 = shift_i_map_30;
      end
      6'b011111 : begin
        _zz_shift_i_1 = shift_i_map_31;
      end
      6'b100000 : begin
        _zz_shift_i_1 = shift_i_map_32;
      end
      6'b100001 : begin
        _zz_shift_i_1 = shift_i_map_33;
      end
      6'b100010 : begin
        _zz_shift_i_1 = shift_i_map_34;
      end
      6'b100011 : begin
        _zz_shift_i_1 = shift_i_map_35;
      end
      6'b100100 : begin
        _zz_shift_i_1 = shift_i_map_36;
      end
      6'b100101 : begin
        _zz_shift_i_1 = shift_i_map_37;
      end
      6'b100110 : begin
        _zz_shift_i_1 = shift_i_map_38;
      end
      default : begin
        _zz_shift_i_1 = shift_i_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_1_1)
      6'b000000 : begin
        _zz_shift_q_1 = shift_q_map_0;
      end
      6'b000001 : begin
        _zz_shift_q_1 = shift_q_map_1;
      end
      6'b000010 : begin
        _zz_shift_q_1 = shift_q_map_2;
      end
      6'b000011 : begin
        _zz_shift_q_1 = shift_q_map_3;
      end
      6'b000100 : begin
        _zz_shift_q_1 = shift_q_map_4;
      end
      6'b000101 : begin
        _zz_shift_q_1 = shift_q_map_5;
      end
      6'b000110 : begin
        _zz_shift_q_1 = shift_q_map_6;
      end
      6'b000111 : begin
        _zz_shift_q_1 = shift_q_map_7;
      end
      6'b001000 : begin
        _zz_shift_q_1 = shift_q_map_8;
      end
      6'b001001 : begin
        _zz_shift_q_1 = shift_q_map_9;
      end
      6'b001010 : begin
        _zz_shift_q_1 = shift_q_map_10;
      end
      6'b001011 : begin
        _zz_shift_q_1 = shift_q_map_11;
      end
      6'b001100 : begin
        _zz_shift_q_1 = shift_q_map_12;
      end
      6'b001101 : begin
        _zz_shift_q_1 = shift_q_map_13;
      end
      6'b001110 : begin
        _zz_shift_q_1 = shift_q_map_14;
      end
      6'b001111 : begin
        _zz_shift_q_1 = shift_q_map_15;
      end
      6'b010000 : begin
        _zz_shift_q_1 = shift_q_map_16;
      end
      6'b010001 : begin
        _zz_shift_q_1 = shift_q_map_17;
      end
      6'b010010 : begin
        _zz_shift_q_1 = shift_q_map_18;
      end
      6'b010011 : begin
        _zz_shift_q_1 = shift_q_map_19;
      end
      6'b010100 : begin
        _zz_shift_q_1 = shift_q_map_20;
      end
      6'b010101 : begin
        _zz_shift_q_1 = shift_q_map_21;
      end
      6'b010110 : begin
        _zz_shift_q_1 = shift_q_map_22;
      end
      6'b010111 : begin
        _zz_shift_q_1 = shift_q_map_23;
      end
      6'b011000 : begin
        _zz_shift_q_1 = shift_q_map_24;
      end
      6'b011001 : begin
        _zz_shift_q_1 = shift_q_map_25;
      end
      6'b011010 : begin
        _zz_shift_q_1 = shift_q_map_26;
      end
      6'b011011 : begin
        _zz_shift_q_1 = shift_q_map_27;
      end
      6'b011100 : begin
        _zz_shift_q_1 = shift_q_map_28;
      end
      6'b011101 : begin
        _zz_shift_q_1 = shift_q_map_29;
      end
      6'b011110 : begin
        _zz_shift_q_1 = shift_q_map_30;
      end
      6'b011111 : begin
        _zz_shift_q_1 = shift_q_map_31;
      end
      6'b100000 : begin
        _zz_shift_q_1 = shift_q_map_32;
      end
      6'b100001 : begin
        _zz_shift_q_1 = shift_q_map_33;
      end
      6'b100010 : begin
        _zz_shift_q_1 = shift_q_map_34;
      end
      6'b100011 : begin
        _zz_shift_q_1 = shift_q_map_35;
      end
      6'b100100 : begin
        _zz_shift_q_1 = shift_q_map_36;
      end
      6'b100101 : begin
        _zz_shift_q_1 = shift_q_map_37;
      end
      6'b100110 : begin
        _zz_shift_q_1 = shift_q_map_38;
      end
      default : begin
        _zz_shift_q_1 = shift_q_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_2_1)
      6'b000000 : begin
        _zz_shift_i_2 = shift_i_map_0;
      end
      6'b000001 : begin
        _zz_shift_i_2 = shift_i_map_1;
      end
      6'b000010 : begin
        _zz_shift_i_2 = shift_i_map_2;
      end
      6'b000011 : begin
        _zz_shift_i_2 = shift_i_map_3;
      end
      6'b000100 : begin
        _zz_shift_i_2 = shift_i_map_4;
      end
      6'b000101 : begin
        _zz_shift_i_2 = shift_i_map_5;
      end
      6'b000110 : begin
        _zz_shift_i_2 = shift_i_map_6;
      end
      6'b000111 : begin
        _zz_shift_i_2 = shift_i_map_7;
      end
      6'b001000 : begin
        _zz_shift_i_2 = shift_i_map_8;
      end
      6'b001001 : begin
        _zz_shift_i_2 = shift_i_map_9;
      end
      6'b001010 : begin
        _zz_shift_i_2 = shift_i_map_10;
      end
      6'b001011 : begin
        _zz_shift_i_2 = shift_i_map_11;
      end
      6'b001100 : begin
        _zz_shift_i_2 = shift_i_map_12;
      end
      6'b001101 : begin
        _zz_shift_i_2 = shift_i_map_13;
      end
      6'b001110 : begin
        _zz_shift_i_2 = shift_i_map_14;
      end
      6'b001111 : begin
        _zz_shift_i_2 = shift_i_map_15;
      end
      6'b010000 : begin
        _zz_shift_i_2 = shift_i_map_16;
      end
      6'b010001 : begin
        _zz_shift_i_2 = shift_i_map_17;
      end
      6'b010010 : begin
        _zz_shift_i_2 = shift_i_map_18;
      end
      6'b010011 : begin
        _zz_shift_i_2 = shift_i_map_19;
      end
      6'b010100 : begin
        _zz_shift_i_2 = shift_i_map_20;
      end
      6'b010101 : begin
        _zz_shift_i_2 = shift_i_map_21;
      end
      6'b010110 : begin
        _zz_shift_i_2 = shift_i_map_22;
      end
      6'b010111 : begin
        _zz_shift_i_2 = shift_i_map_23;
      end
      6'b011000 : begin
        _zz_shift_i_2 = shift_i_map_24;
      end
      6'b011001 : begin
        _zz_shift_i_2 = shift_i_map_25;
      end
      6'b011010 : begin
        _zz_shift_i_2 = shift_i_map_26;
      end
      6'b011011 : begin
        _zz_shift_i_2 = shift_i_map_27;
      end
      6'b011100 : begin
        _zz_shift_i_2 = shift_i_map_28;
      end
      6'b011101 : begin
        _zz_shift_i_2 = shift_i_map_29;
      end
      6'b011110 : begin
        _zz_shift_i_2 = shift_i_map_30;
      end
      6'b011111 : begin
        _zz_shift_i_2 = shift_i_map_31;
      end
      6'b100000 : begin
        _zz_shift_i_2 = shift_i_map_32;
      end
      6'b100001 : begin
        _zz_shift_i_2 = shift_i_map_33;
      end
      6'b100010 : begin
        _zz_shift_i_2 = shift_i_map_34;
      end
      6'b100011 : begin
        _zz_shift_i_2 = shift_i_map_35;
      end
      6'b100100 : begin
        _zz_shift_i_2 = shift_i_map_36;
      end
      6'b100101 : begin
        _zz_shift_i_2 = shift_i_map_37;
      end
      6'b100110 : begin
        _zz_shift_i_2 = shift_i_map_38;
      end
      default : begin
        _zz_shift_i_2 = shift_i_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_2_1)
      6'b000000 : begin
        _zz_shift_q_2 = shift_q_map_0;
      end
      6'b000001 : begin
        _zz_shift_q_2 = shift_q_map_1;
      end
      6'b000010 : begin
        _zz_shift_q_2 = shift_q_map_2;
      end
      6'b000011 : begin
        _zz_shift_q_2 = shift_q_map_3;
      end
      6'b000100 : begin
        _zz_shift_q_2 = shift_q_map_4;
      end
      6'b000101 : begin
        _zz_shift_q_2 = shift_q_map_5;
      end
      6'b000110 : begin
        _zz_shift_q_2 = shift_q_map_6;
      end
      6'b000111 : begin
        _zz_shift_q_2 = shift_q_map_7;
      end
      6'b001000 : begin
        _zz_shift_q_2 = shift_q_map_8;
      end
      6'b001001 : begin
        _zz_shift_q_2 = shift_q_map_9;
      end
      6'b001010 : begin
        _zz_shift_q_2 = shift_q_map_10;
      end
      6'b001011 : begin
        _zz_shift_q_2 = shift_q_map_11;
      end
      6'b001100 : begin
        _zz_shift_q_2 = shift_q_map_12;
      end
      6'b001101 : begin
        _zz_shift_q_2 = shift_q_map_13;
      end
      6'b001110 : begin
        _zz_shift_q_2 = shift_q_map_14;
      end
      6'b001111 : begin
        _zz_shift_q_2 = shift_q_map_15;
      end
      6'b010000 : begin
        _zz_shift_q_2 = shift_q_map_16;
      end
      6'b010001 : begin
        _zz_shift_q_2 = shift_q_map_17;
      end
      6'b010010 : begin
        _zz_shift_q_2 = shift_q_map_18;
      end
      6'b010011 : begin
        _zz_shift_q_2 = shift_q_map_19;
      end
      6'b010100 : begin
        _zz_shift_q_2 = shift_q_map_20;
      end
      6'b010101 : begin
        _zz_shift_q_2 = shift_q_map_21;
      end
      6'b010110 : begin
        _zz_shift_q_2 = shift_q_map_22;
      end
      6'b010111 : begin
        _zz_shift_q_2 = shift_q_map_23;
      end
      6'b011000 : begin
        _zz_shift_q_2 = shift_q_map_24;
      end
      6'b011001 : begin
        _zz_shift_q_2 = shift_q_map_25;
      end
      6'b011010 : begin
        _zz_shift_q_2 = shift_q_map_26;
      end
      6'b011011 : begin
        _zz_shift_q_2 = shift_q_map_27;
      end
      6'b011100 : begin
        _zz_shift_q_2 = shift_q_map_28;
      end
      6'b011101 : begin
        _zz_shift_q_2 = shift_q_map_29;
      end
      6'b011110 : begin
        _zz_shift_q_2 = shift_q_map_30;
      end
      6'b011111 : begin
        _zz_shift_q_2 = shift_q_map_31;
      end
      6'b100000 : begin
        _zz_shift_q_2 = shift_q_map_32;
      end
      6'b100001 : begin
        _zz_shift_q_2 = shift_q_map_33;
      end
      6'b100010 : begin
        _zz_shift_q_2 = shift_q_map_34;
      end
      6'b100011 : begin
        _zz_shift_q_2 = shift_q_map_35;
      end
      6'b100100 : begin
        _zz_shift_q_2 = shift_q_map_36;
      end
      6'b100101 : begin
        _zz_shift_q_2 = shift_q_map_37;
      end
      6'b100110 : begin
        _zz_shift_q_2 = shift_q_map_38;
      end
      default : begin
        _zz_shift_q_2 = shift_q_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_3_1)
      6'b000000 : begin
        _zz_shift_i_3 = shift_i_map_0;
      end
      6'b000001 : begin
        _zz_shift_i_3 = shift_i_map_1;
      end
      6'b000010 : begin
        _zz_shift_i_3 = shift_i_map_2;
      end
      6'b000011 : begin
        _zz_shift_i_3 = shift_i_map_3;
      end
      6'b000100 : begin
        _zz_shift_i_3 = shift_i_map_4;
      end
      6'b000101 : begin
        _zz_shift_i_3 = shift_i_map_5;
      end
      6'b000110 : begin
        _zz_shift_i_3 = shift_i_map_6;
      end
      6'b000111 : begin
        _zz_shift_i_3 = shift_i_map_7;
      end
      6'b001000 : begin
        _zz_shift_i_3 = shift_i_map_8;
      end
      6'b001001 : begin
        _zz_shift_i_3 = shift_i_map_9;
      end
      6'b001010 : begin
        _zz_shift_i_3 = shift_i_map_10;
      end
      6'b001011 : begin
        _zz_shift_i_3 = shift_i_map_11;
      end
      6'b001100 : begin
        _zz_shift_i_3 = shift_i_map_12;
      end
      6'b001101 : begin
        _zz_shift_i_3 = shift_i_map_13;
      end
      6'b001110 : begin
        _zz_shift_i_3 = shift_i_map_14;
      end
      6'b001111 : begin
        _zz_shift_i_3 = shift_i_map_15;
      end
      6'b010000 : begin
        _zz_shift_i_3 = shift_i_map_16;
      end
      6'b010001 : begin
        _zz_shift_i_3 = shift_i_map_17;
      end
      6'b010010 : begin
        _zz_shift_i_3 = shift_i_map_18;
      end
      6'b010011 : begin
        _zz_shift_i_3 = shift_i_map_19;
      end
      6'b010100 : begin
        _zz_shift_i_3 = shift_i_map_20;
      end
      6'b010101 : begin
        _zz_shift_i_3 = shift_i_map_21;
      end
      6'b010110 : begin
        _zz_shift_i_3 = shift_i_map_22;
      end
      6'b010111 : begin
        _zz_shift_i_3 = shift_i_map_23;
      end
      6'b011000 : begin
        _zz_shift_i_3 = shift_i_map_24;
      end
      6'b011001 : begin
        _zz_shift_i_3 = shift_i_map_25;
      end
      6'b011010 : begin
        _zz_shift_i_3 = shift_i_map_26;
      end
      6'b011011 : begin
        _zz_shift_i_3 = shift_i_map_27;
      end
      6'b011100 : begin
        _zz_shift_i_3 = shift_i_map_28;
      end
      6'b011101 : begin
        _zz_shift_i_3 = shift_i_map_29;
      end
      6'b011110 : begin
        _zz_shift_i_3 = shift_i_map_30;
      end
      6'b011111 : begin
        _zz_shift_i_3 = shift_i_map_31;
      end
      6'b100000 : begin
        _zz_shift_i_3 = shift_i_map_32;
      end
      6'b100001 : begin
        _zz_shift_i_3 = shift_i_map_33;
      end
      6'b100010 : begin
        _zz_shift_i_3 = shift_i_map_34;
      end
      6'b100011 : begin
        _zz_shift_i_3 = shift_i_map_35;
      end
      6'b100100 : begin
        _zz_shift_i_3 = shift_i_map_36;
      end
      6'b100101 : begin
        _zz_shift_i_3 = shift_i_map_37;
      end
      6'b100110 : begin
        _zz_shift_i_3 = shift_i_map_38;
      end
      default : begin
        _zz_shift_i_3 = shift_i_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_3_1)
      6'b000000 : begin
        _zz_shift_q_3 = shift_q_map_0;
      end
      6'b000001 : begin
        _zz_shift_q_3 = shift_q_map_1;
      end
      6'b000010 : begin
        _zz_shift_q_3 = shift_q_map_2;
      end
      6'b000011 : begin
        _zz_shift_q_3 = shift_q_map_3;
      end
      6'b000100 : begin
        _zz_shift_q_3 = shift_q_map_4;
      end
      6'b000101 : begin
        _zz_shift_q_3 = shift_q_map_5;
      end
      6'b000110 : begin
        _zz_shift_q_3 = shift_q_map_6;
      end
      6'b000111 : begin
        _zz_shift_q_3 = shift_q_map_7;
      end
      6'b001000 : begin
        _zz_shift_q_3 = shift_q_map_8;
      end
      6'b001001 : begin
        _zz_shift_q_3 = shift_q_map_9;
      end
      6'b001010 : begin
        _zz_shift_q_3 = shift_q_map_10;
      end
      6'b001011 : begin
        _zz_shift_q_3 = shift_q_map_11;
      end
      6'b001100 : begin
        _zz_shift_q_3 = shift_q_map_12;
      end
      6'b001101 : begin
        _zz_shift_q_3 = shift_q_map_13;
      end
      6'b001110 : begin
        _zz_shift_q_3 = shift_q_map_14;
      end
      6'b001111 : begin
        _zz_shift_q_3 = shift_q_map_15;
      end
      6'b010000 : begin
        _zz_shift_q_3 = shift_q_map_16;
      end
      6'b010001 : begin
        _zz_shift_q_3 = shift_q_map_17;
      end
      6'b010010 : begin
        _zz_shift_q_3 = shift_q_map_18;
      end
      6'b010011 : begin
        _zz_shift_q_3 = shift_q_map_19;
      end
      6'b010100 : begin
        _zz_shift_q_3 = shift_q_map_20;
      end
      6'b010101 : begin
        _zz_shift_q_3 = shift_q_map_21;
      end
      6'b010110 : begin
        _zz_shift_q_3 = shift_q_map_22;
      end
      6'b010111 : begin
        _zz_shift_q_3 = shift_q_map_23;
      end
      6'b011000 : begin
        _zz_shift_q_3 = shift_q_map_24;
      end
      6'b011001 : begin
        _zz_shift_q_3 = shift_q_map_25;
      end
      6'b011010 : begin
        _zz_shift_q_3 = shift_q_map_26;
      end
      6'b011011 : begin
        _zz_shift_q_3 = shift_q_map_27;
      end
      6'b011100 : begin
        _zz_shift_q_3 = shift_q_map_28;
      end
      6'b011101 : begin
        _zz_shift_q_3 = shift_q_map_29;
      end
      6'b011110 : begin
        _zz_shift_q_3 = shift_q_map_30;
      end
      6'b011111 : begin
        _zz_shift_q_3 = shift_q_map_31;
      end
      6'b100000 : begin
        _zz_shift_q_3 = shift_q_map_32;
      end
      6'b100001 : begin
        _zz_shift_q_3 = shift_q_map_33;
      end
      6'b100010 : begin
        _zz_shift_q_3 = shift_q_map_34;
      end
      6'b100011 : begin
        _zz_shift_q_3 = shift_q_map_35;
      end
      6'b100100 : begin
        _zz_shift_q_3 = shift_q_map_36;
      end
      6'b100101 : begin
        _zz_shift_q_3 = shift_q_map_37;
      end
      6'b100110 : begin
        _zz_shift_q_3 = shift_q_map_38;
      end
      default : begin
        _zz_shift_q_3 = shift_q_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_4_1)
      6'b000000 : begin
        _zz_shift_i_4 = shift_i_map_0;
      end
      6'b000001 : begin
        _zz_shift_i_4 = shift_i_map_1;
      end
      6'b000010 : begin
        _zz_shift_i_4 = shift_i_map_2;
      end
      6'b000011 : begin
        _zz_shift_i_4 = shift_i_map_3;
      end
      6'b000100 : begin
        _zz_shift_i_4 = shift_i_map_4;
      end
      6'b000101 : begin
        _zz_shift_i_4 = shift_i_map_5;
      end
      6'b000110 : begin
        _zz_shift_i_4 = shift_i_map_6;
      end
      6'b000111 : begin
        _zz_shift_i_4 = shift_i_map_7;
      end
      6'b001000 : begin
        _zz_shift_i_4 = shift_i_map_8;
      end
      6'b001001 : begin
        _zz_shift_i_4 = shift_i_map_9;
      end
      6'b001010 : begin
        _zz_shift_i_4 = shift_i_map_10;
      end
      6'b001011 : begin
        _zz_shift_i_4 = shift_i_map_11;
      end
      6'b001100 : begin
        _zz_shift_i_4 = shift_i_map_12;
      end
      6'b001101 : begin
        _zz_shift_i_4 = shift_i_map_13;
      end
      6'b001110 : begin
        _zz_shift_i_4 = shift_i_map_14;
      end
      6'b001111 : begin
        _zz_shift_i_4 = shift_i_map_15;
      end
      6'b010000 : begin
        _zz_shift_i_4 = shift_i_map_16;
      end
      6'b010001 : begin
        _zz_shift_i_4 = shift_i_map_17;
      end
      6'b010010 : begin
        _zz_shift_i_4 = shift_i_map_18;
      end
      6'b010011 : begin
        _zz_shift_i_4 = shift_i_map_19;
      end
      6'b010100 : begin
        _zz_shift_i_4 = shift_i_map_20;
      end
      6'b010101 : begin
        _zz_shift_i_4 = shift_i_map_21;
      end
      6'b010110 : begin
        _zz_shift_i_4 = shift_i_map_22;
      end
      6'b010111 : begin
        _zz_shift_i_4 = shift_i_map_23;
      end
      6'b011000 : begin
        _zz_shift_i_4 = shift_i_map_24;
      end
      6'b011001 : begin
        _zz_shift_i_4 = shift_i_map_25;
      end
      6'b011010 : begin
        _zz_shift_i_4 = shift_i_map_26;
      end
      6'b011011 : begin
        _zz_shift_i_4 = shift_i_map_27;
      end
      6'b011100 : begin
        _zz_shift_i_4 = shift_i_map_28;
      end
      6'b011101 : begin
        _zz_shift_i_4 = shift_i_map_29;
      end
      6'b011110 : begin
        _zz_shift_i_4 = shift_i_map_30;
      end
      6'b011111 : begin
        _zz_shift_i_4 = shift_i_map_31;
      end
      6'b100000 : begin
        _zz_shift_i_4 = shift_i_map_32;
      end
      6'b100001 : begin
        _zz_shift_i_4 = shift_i_map_33;
      end
      6'b100010 : begin
        _zz_shift_i_4 = shift_i_map_34;
      end
      6'b100011 : begin
        _zz_shift_i_4 = shift_i_map_35;
      end
      6'b100100 : begin
        _zz_shift_i_4 = shift_i_map_36;
      end
      6'b100101 : begin
        _zz_shift_i_4 = shift_i_map_37;
      end
      6'b100110 : begin
        _zz_shift_i_4 = shift_i_map_38;
      end
      default : begin
        _zz_shift_i_4 = shift_i_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_4_1)
      6'b000000 : begin
        _zz_shift_q_4 = shift_q_map_0;
      end
      6'b000001 : begin
        _zz_shift_q_4 = shift_q_map_1;
      end
      6'b000010 : begin
        _zz_shift_q_4 = shift_q_map_2;
      end
      6'b000011 : begin
        _zz_shift_q_4 = shift_q_map_3;
      end
      6'b000100 : begin
        _zz_shift_q_4 = shift_q_map_4;
      end
      6'b000101 : begin
        _zz_shift_q_4 = shift_q_map_5;
      end
      6'b000110 : begin
        _zz_shift_q_4 = shift_q_map_6;
      end
      6'b000111 : begin
        _zz_shift_q_4 = shift_q_map_7;
      end
      6'b001000 : begin
        _zz_shift_q_4 = shift_q_map_8;
      end
      6'b001001 : begin
        _zz_shift_q_4 = shift_q_map_9;
      end
      6'b001010 : begin
        _zz_shift_q_4 = shift_q_map_10;
      end
      6'b001011 : begin
        _zz_shift_q_4 = shift_q_map_11;
      end
      6'b001100 : begin
        _zz_shift_q_4 = shift_q_map_12;
      end
      6'b001101 : begin
        _zz_shift_q_4 = shift_q_map_13;
      end
      6'b001110 : begin
        _zz_shift_q_4 = shift_q_map_14;
      end
      6'b001111 : begin
        _zz_shift_q_4 = shift_q_map_15;
      end
      6'b010000 : begin
        _zz_shift_q_4 = shift_q_map_16;
      end
      6'b010001 : begin
        _zz_shift_q_4 = shift_q_map_17;
      end
      6'b010010 : begin
        _zz_shift_q_4 = shift_q_map_18;
      end
      6'b010011 : begin
        _zz_shift_q_4 = shift_q_map_19;
      end
      6'b010100 : begin
        _zz_shift_q_4 = shift_q_map_20;
      end
      6'b010101 : begin
        _zz_shift_q_4 = shift_q_map_21;
      end
      6'b010110 : begin
        _zz_shift_q_4 = shift_q_map_22;
      end
      6'b010111 : begin
        _zz_shift_q_4 = shift_q_map_23;
      end
      6'b011000 : begin
        _zz_shift_q_4 = shift_q_map_24;
      end
      6'b011001 : begin
        _zz_shift_q_4 = shift_q_map_25;
      end
      6'b011010 : begin
        _zz_shift_q_4 = shift_q_map_26;
      end
      6'b011011 : begin
        _zz_shift_q_4 = shift_q_map_27;
      end
      6'b011100 : begin
        _zz_shift_q_4 = shift_q_map_28;
      end
      6'b011101 : begin
        _zz_shift_q_4 = shift_q_map_29;
      end
      6'b011110 : begin
        _zz_shift_q_4 = shift_q_map_30;
      end
      6'b011111 : begin
        _zz_shift_q_4 = shift_q_map_31;
      end
      6'b100000 : begin
        _zz_shift_q_4 = shift_q_map_32;
      end
      6'b100001 : begin
        _zz_shift_q_4 = shift_q_map_33;
      end
      6'b100010 : begin
        _zz_shift_q_4 = shift_q_map_34;
      end
      6'b100011 : begin
        _zz_shift_q_4 = shift_q_map_35;
      end
      6'b100100 : begin
        _zz_shift_q_4 = shift_q_map_36;
      end
      6'b100101 : begin
        _zz_shift_q_4 = shift_q_map_37;
      end
      6'b100110 : begin
        _zz_shift_q_4 = shift_q_map_38;
      end
      default : begin
        _zz_shift_q_4 = shift_q_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_5_1)
      6'b000000 : begin
        _zz_shift_i_5 = shift_i_map_0;
      end
      6'b000001 : begin
        _zz_shift_i_5 = shift_i_map_1;
      end
      6'b000010 : begin
        _zz_shift_i_5 = shift_i_map_2;
      end
      6'b000011 : begin
        _zz_shift_i_5 = shift_i_map_3;
      end
      6'b000100 : begin
        _zz_shift_i_5 = shift_i_map_4;
      end
      6'b000101 : begin
        _zz_shift_i_5 = shift_i_map_5;
      end
      6'b000110 : begin
        _zz_shift_i_5 = shift_i_map_6;
      end
      6'b000111 : begin
        _zz_shift_i_5 = shift_i_map_7;
      end
      6'b001000 : begin
        _zz_shift_i_5 = shift_i_map_8;
      end
      6'b001001 : begin
        _zz_shift_i_5 = shift_i_map_9;
      end
      6'b001010 : begin
        _zz_shift_i_5 = shift_i_map_10;
      end
      6'b001011 : begin
        _zz_shift_i_5 = shift_i_map_11;
      end
      6'b001100 : begin
        _zz_shift_i_5 = shift_i_map_12;
      end
      6'b001101 : begin
        _zz_shift_i_5 = shift_i_map_13;
      end
      6'b001110 : begin
        _zz_shift_i_5 = shift_i_map_14;
      end
      6'b001111 : begin
        _zz_shift_i_5 = shift_i_map_15;
      end
      6'b010000 : begin
        _zz_shift_i_5 = shift_i_map_16;
      end
      6'b010001 : begin
        _zz_shift_i_5 = shift_i_map_17;
      end
      6'b010010 : begin
        _zz_shift_i_5 = shift_i_map_18;
      end
      6'b010011 : begin
        _zz_shift_i_5 = shift_i_map_19;
      end
      6'b010100 : begin
        _zz_shift_i_5 = shift_i_map_20;
      end
      6'b010101 : begin
        _zz_shift_i_5 = shift_i_map_21;
      end
      6'b010110 : begin
        _zz_shift_i_5 = shift_i_map_22;
      end
      6'b010111 : begin
        _zz_shift_i_5 = shift_i_map_23;
      end
      6'b011000 : begin
        _zz_shift_i_5 = shift_i_map_24;
      end
      6'b011001 : begin
        _zz_shift_i_5 = shift_i_map_25;
      end
      6'b011010 : begin
        _zz_shift_i_5 = shift_i_map_26;
      end
      6'b011011 : begin
        _zz_shift_i_5 = shift_i_map_27;
      end
      6'b011100 : begin
        _zz_shift_i_5 = shift_i_map_28;
      end
      6'b011101 : begin
        _zz_shift_i_5 = shift_i_map_29;
      end
      6'b011110 : begin
        _zz_shift_i_5 = shift_i_map_30;
      end
      6'b011111 : begin
        _zz_shift_i_5 = shift_i_map_31;
      end
      6'b100000 : begin
        _zz_shift_i_5 = shift_i_map_32;
      end
      6'b100001 : begin
        _zz_shift_i_5 = shift_i_map_33;
      end
      6'b100010 : begin
        _zz_shift_i_5 = shift_i_map_34;
      end
      6'b100011 : begin
        _zz_shift_i_5 = shift_i_map_35;
      end
      6'b100100 : begin
        _zz_shift_i_5 = shift_i_map_36;
      end
      6'b100101 : begin
        _zz_shift_i_5 = shift_i_map_37;
      end
      6'b100110 : begin
        _zz_shift_i_5 = shift_i_map_38;
      end
      default : begin
        _zz_shift_i_5 = shift_i_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_5_1)
      6'b000000 : begin
        _zz_shift_q_5 = shift_q_map_0;
      end
      6'b000001 : begin
        _zz_shift_q_5 = shift_q_map_1;
      end
      6'b000010 : begin
        _zz_shift_q_5 = shift_q_map_2;
      end
      6'b000011 : begin
        _zz_shift_q_5 = shift_q_map_3;
      end
      6'b000100 : begin
        _zz_shift_q_5 = shift_q_map_4;
      end
      6'b000101 : begin
        _zz_shift_q_5 = shift_q_map_5;
      end
      6'b000110 : begin
        _zz_shift_q_5 = shift_q_map_6;
      end
      6'b000111 : begin
        _zz_shift_q_5 = shift_q_map_7;
      end
      6'b001000 : begin
        _zz_shift_q_5 = shift_q_map_8;
      end
      6'b001001 : begin
        _zz_shift_q_5 = shift_q_map_9;
      end
      6'b001010 : begin
        _zz_shift_q_5 = shift_q_map_10;
      end
      6'b001011 : begin
        _zz_shift_q_5 = shift_q_map_11;
      end
      6'b001100 : begin
        _zz_shift_q_5 = shift_q_map_12;
      end
      6'b001101 : begin
        _zz_shift_q_5 = shift_q_map_13;
      end
      6'b001110 : begin
        _zz_shift_q_5 = shift_q_map_14;
      end
      6'b001111 : begin
        _zz_shift_q_5 = shift_q_map_15;
      end
      6'b010000 : begin
        _zz_shift_q_5 = shift_q_map_16;
      end
      6'b010001 : begin
        _zz_shift_q_5 = shift_q_map_17;
      end
      6'b010010 : begin
        _zz_shift_q_5 = shift_q_map_18;
      end
      6'b010011 : begin
        _zz_shift_q_5 = shift_q_map_19;
      end
      6'b010100 : begin
        _zz_shift_q_5 = shift_q_map_20;
      end
      6'b010101 : begin
        _zz_shift_q_5 = shift_q_map_21;
      end
      6'b010110 : begin
        _zz_shift_q_5 = shift_q_map_22;
      end
      6'b010111 : begin
        _zz_shift_q_5 = shift_q_map_23;
      end
      6'b011000 : begin
        _zz_shift_q_5 = shift_q_map_24;
      end
      6'b011001 : begin
        _zz_shift_q_5 = shift_q_map_25;
      end
      6'b011010 : begin
        _zz_shift_q_5 = shift_q_map_26;
      end
      6'b011011 : begin
        _zz_shift_q_5 = shift_q_map_27;
      end
      6'b011100 : begin
        _zz_shift_q_5 = shift_q_map_28;
      end
      6'b011101 : begin
        _zz_shift_q_5 = shift_q_map_29;
      end
      6'b011110 : begin
        _zz_shift_q_5 = shift_q_map_30;
      end
      6'b011111 : begin
        _zz_shift_q_5 = shift_q_map_31;
      end
      6'b100000 : begin
        _zz_shift_q_5 = shift_q_map_32;
      end
      6'b100001 : begin
        _zz_shift_q_5 = shift_q_map_33;
      end
      6'b100010 : begin
        _zz_shift_q_5 = shift_q_map_34;
      end
      6'b100011 : begin
        _zz_shift_q_5 = shift_q_map_35;
      end
      6'b100100 : begin
        _zz_shift_q_5 = shift_q_map_36;
      end
      6'b100101 : begin
        _zz_shift_q_5 = shift_q_map_37;
      end
      6'b100110 : begin
        _zz_shift_q_5 = shift_q_map_38;
      end
      default : begin
        _zz_shift_q_5 = shift_q_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_6_1)
      6'b000000 : begin
        _zz_shift_i_6 = shift_i_map_0;
      end
      6'b000001 : begin
        _zz_shift_i_6 = shift_i_map_1;
      end
      6'b000010 : begin
        _zz_shift_i_6 = shift_i_map_2;
      end
      6'b000011 : begin
        _zz_shift_i_6 = shift_i_map_3;
      end
      6'b000100 : begin
        _zz_shift_i_6 = shift_i_map_4;
      end
      6'b000101 : begin
        _zz_shift_i_6 = shift_i_map_5;
      end
      6'b000110 : begin
        _zz_shift_i_6 = shift_i_map_6;
      end
      6'b000111 : begin
        _zz_shift_i_6 = shift_i_map_7;
      end
      6'b001000 : begin
        _zz_shift_i_6 = shift_i_map_8;
      end
      6'b001001 : begin
        _zz_shift_i_6 = shift_i_map_9;
      end
      6'b001010 : begin
        _zz_shift_i_6 = shift_i_map_10;
      end
      6'b001011 : begin
        _zz_shift_i_6 = shift_i_map_11;
      end
      6'b001100 : begin
        _zz_shift_i_6 = shift_i_map_12;
      end
      6'b001101 : begin
        _zz_shift_i_6 = shift_i_map_13;
      end
      6'b001110 : begin
        _zz_shift_i_6 = shift_i_map_14;
      end
      6'b001111 : begin
        _zz_shift_i_6 = shift_i_map_15;
      end
      6'b010000 : begin
        _zz_shift_i_6 = shift_i_map_16;
      end
      6'b010001 : begin
        _zz_shift_i_6 = shift_i_map_17;
      end
      6'b010010 : begin
        _zz_shift_i_6 = shift_i_map_18;
      end
      6'b010011 : begin
        _zz_shift_i_6 = shift_i_map_19;
      end
      6'b010100 : begin
        _zz_shift_i_6 = shift_i_map_20;
      end
      6'b010101 : begin
        _zz_shift_i_6 = shift_i_map_21;
      end
      6'b010110 : begin
        _zz_shift_i_6 = shift_i_map_22;
      end
      6'b010111 : begin
        _zz_shift_i_6 = shift_i_map_23;
      end
      6'b011000 : begin
        _zz_shift_i_6 = shift_i_map_24;
      end
      6'b011001 : begin
        _zz_shift_i_6 = shift_i_map_25;
      end
      6'b011010 : begin
        _zz_shift_i_6 = shift_i_map_26;
      end
      6'b011011 : begin
        _zz_shift_i_6 = shift_i_map_27;
      end
      6'b011100 : begin
        _zz_shift_i_6 = shift_i_map_28;
      end
      6'b011101 : begin
        _zz_shift_i_6 = shift_i_map_29;
      end
      6'b011110 : begin
        _zz_shift_i_6 = shift_i_map_30;
      end
      6'b011111 : begin
        _zz_shift_i_6 = shift_i_map_31;
      end
      6'b100000 : begin
        _zz_shift_i_6 = shift_i_map_32;
      end
      6'b100001 : begin
        _zz_shift_i_6 = shift_i_map_33;
      end
      6'b100010 : begin
        _zz_shift_i_6 = shift_i_map_34;
      end
      6'b100011 : begin
        _zz_shift_i_6 = shift_i_map_35;
      end
      6'b100100 : begin
        _zz_shift_i_6 = shift_i_map_36;
      end
      6'b100101 : begin
        _zz_shift_i_6 = shift_i_map_37;
      end
      6'b100110 : begin
        _zz_shift_i_6 = shift_i_map_38;
      end
      default : begin
        _zz_shift_i_6 = shift_i_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_6_1)
      6'b000000 : begin
        _zz_shift_q_6 = shift_q_map_0;
      end
      6'b000001 : begin
        _zz_shift_q_6 = shift_q_map_1;
      end
      6'b000010 : begin
        _zz_shift_q_6 = shift_q_map_2;
      end
      6'b000011 : begin
        _zz_shift_q_6 = shift_q_map_3;
      end
      6'b000100 : begin
        _zz_shift_q_6 = shift_q_map_4;
      end
      6'b000101 : begin
        _zz_shift_q_6 = shift_q_map_5;
      end
      6'b000110 : begin
        _zz_shift_q_6 = shift_q_map_6;
      end
      6'b000111 : begin
        _zz_shift_q_6 = shift_q_map_7;
      end
      6'b001000 : begin
        _zz_shift_q_6 = shift_q_map_8;
      end
      6'b001001 : begin
        _zz_shift_q_6 = shift_q_map_9;
      end
      6'b001010 : begin
        _zz_shift_q_6 = shift_q_map_10;
      end
      6'b001011 : begin
        _zz_shift_q_6 = shift_q_map_11;
      end
      6'b001100 : begin
        _zz_shift_q_6 = shift_q_map_12;
      end
      6'b001101 : begin
        _zz_shift_q_6 = shift_q_map_13;
      end
      6'b001110 : begin
        _zz_shift_q_6 = shift_q_map_14;
      end
      6'b001111 : begin
        _zz_shift_q_6 = shift_q_map_15;
      end
      6'b010000 : begin
        _zz_shift_q_6 = shift_q_map_16;
      end
      6'b010001 : begin
        _zz_shift_q_6 = shift_q_map_17;
      end
      6'b010010 : begin
        _zz_shift_q_6 = shift_q_map_18;
      end
      6'b010011 : begin
        _zz_shift_q_6 = shift_q_map_19;
      end
      6'b010100 : begin
        _zz_shift_q_6 = shift_q_map_20;
      end
      6'b010101 : begin
        _zz_shift_q_6 = shift_q_map_21;
      end
      6'b010110 : begin
        _zz_shift_q_6 = shift_q_map_22;
      end
      6'b010111 : begin
        _zz_shift_q_6 = shift_q_map_23;
      end
      6'b011000 : begin
        _zz_shift_q_6 = shift_q_map_24;
      end
      6'b011001 : begin
        _zz_shift_q_6 = shift_q_map_25;
      end
      6'b011010 : begin
        _zz_shift_q_6 = shift_q_map_26;
      end
      6'b011011 : begin
        _zz_shift_q_6 = shift_q_map_27;
      end
      6'b011100 : begin
        _zz_shift_q_6 = shift_q_map_28;
      end
      6'b011101 : begin
        _zz_shift_q_6 = shift_q_map_29;
      end
      6'b011110 : begin
        _zz_shift_q_6 = shift_q_map_30;
      end
      6'b011111 : begin
        _zz_shift_q_6 = shift_q_map_31;
      end
      6'b100000 : begin
        _zz_shift_q_6 = shift_q_map_32;
      end
      6'b100001 : begin
        _zz_shift_q_6 = shift_q_map_33;
      end
      6'b100010 : begin
        _zz_shift_q_6 = shift_q_map_34;
      end
      6'b100011 : begin
        _zz_shift_q_6 = shift_q_map_35;
      end
      6'b100100 : begin
        _zz_shift_q_6 = shift_q_map_36;
      end
      6'b100101 : begin
        _zz_shift_q_6 = shift_q_map_37;
      end
      6'b100110 : begin
        _zz_shift_q_6 = shift_q_map_38;
      end
      default : begin
        _zz_shift_q_6 = shift_q_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_7_1)
      6'b000000 : begin
        _zz_shift_i_7 = shift_i_map_0;
      end
      6'b000001 : begin
        _zz_shift_i_7 = shift_i_map_1;
      end
      6'b000010 : begin
        _zz_shift_i_7 = shift_i_map_2;
      end
      6'b000011 : begin
        _zz_shift_i_7 = shift_i_map_3;
      end
      6'b000100 : begin
        _zz_shift_i_7 = shift_i_map_4;
      end
      6'b000101 : begin
        _zz_shift_i_7 = shift_i_map_5;
      end
      6'b000110 : begin
        _zz_shift_i_7 = shift_i_map_6;
      end
      6'b000111 : begin
        _zz_shift_i_7 = shift_i_map_7;
      end
      6'b001000 : begin
        _zz_shift_i_7 = shift_i_map_8;
      end
      6'b001001 : begin
        _zz_shift_i_7 = shift_i_map_9;
      end
      6'b001010 : begin
        _zz_shift_i_7 = shift_i_map_10;
      end
      6'b001011 : begin
        _zz_shift_i_7 = shift_i_map_11;
      end
      6'b001100 : begin
        _zz_shift_i_7 = shift_i_map_12;
      end
      6'b001101 : begin
        _zz_shift_i_7 = shift_i_map_13;
      end
      6'b001110 : begin
        _zz_shift_i_7 = shift_i_map_14;
      end
      6'b001111 : begin
        _zz_shift_i_7 = shift_i_map_15;
      end
      6'b010000 : begin
        _zz_shift_i_7 = shift_i_map_16;
      end
      6'b010001 : begin
        _zz_shift_i_7 = shift_i_map_17;
      end
      6'b010010 : begin
        _zz_shift_i_7 = shift_i_map_18;
      end
      6'b010011 : begin
        _zz_shift_i_7 = shift_i_map_19;
      end
      6'b010100 : begin
        _zz_shift_i_7 = shift_i_map_20;
      end
      6'b010101 : begin
        _zz_shift_i_7 = shift_i_map_21;
      end
      6'b010110 : begin
        _zz_shift_i_7 = shift_i_map_22;
      end
      6'b010111 : begin
        _zz_shift_i_7 = shift_i_map_23;
      end
      6'b011000 : begin
        _zz_shift_i_7 = shift_i_map_24;
      end
      6'b011001 : begin
        _zz_shift_i_7 = shift_i_map_25;
      end
      6'b011010 : begin
        _zz_shift_i_7 = shift_i_map_26;
      end
      6'b011011 : begin
        _zz_shift_i_7 = shift_i_map_27;
      end
      6'b011100 : begin
        _zz_shift_i_7 = shift_i_map_28;
      end
      6'b011101 : begin
        _zz_shift_i_7 = shift_i_map_29;
      end
      6'b011110 : begin
        _zz_shift_i_7 = shift_i_map_30;
      end
      6'b011111 : begin
        _zz_shift_i_7 = shift_i_map_31;
      end
      6'b100000 : begin
        _zz_shift_i_7 = shift_i_map_32;
      end
      6'b100001 : begin
        _zz_shift_i_7 = shift_i_map_33;
      end
      6'b100010 : begin
        _zz_shift_i_7 = shift_i_map_34;
      end
      6'b100011 : begin
        _zz_shift_i_7 = shift_i_map_35;
      end
      6'b100100 : begin
        _zz_shift_i_7 = shift_i_map_36;
      end
      6'b100101 : begin
        _zz_shift_i_7 = shift_i_map_37;
      end
      6'b100110 : begin
        _zz_shift_i_7 = shift_i_map_38;
      end
      default : begin
        _zz_shift_i_7 = shift_i_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_7_1)
      6'b000000 : begin
        _zz_shift_q_7 = shift_q_map_0;
      end
      6'b000001 : begin
        _zz_shift_q_7 = shift_q_map_1;
      end
      6'b000010 : begin
        _zz_shift_q_7 = shift_q_map_2;
      end
      6'b000011 : begin
        _zz_shift_q_7 = shift_q_map_3;
      end
      6'b000100 : begin
        _zz_shift_q_7 = shift_q_map_4;
      end
      6'b000101 : begin
        _zz_shift_q_7 = shift_q_map_5;
      end
      6'b000110 : begin
        _zz_shift_q_7 = shift_q_map_6;
      end
      6'b000111 : begin
        _zz_shift_q_7 = shift_q_map_7;
      end
      6'b001000 : begin
        _zz_shift_q_7 = shift_q_map_8;
      end
      6'b001001 : begin
        _zz_shift_q_7 = shift_q_map_9;
      end
      6'b001010 : begin
        _zz_shift_q_7 = shift_q_map_10;
      end
      6'b001011 : begin
        _zz_shift_q_7 = shift_q_map_11;
      end
      6'b001100 : begin
        _zz_shift_q_7 = shift_q_map_12;
      end
      6'b001101 : begin
        _zz_shift_q_7 = shift_q_map_13;
      end
      6'b001110 : begin
        _zz_shift_q_7 = shift_q_map_14;
      end
      6'b001111 : begin
        _zz_shift_q_7 = shift_q_map_15;
      end
      6'b010000 : begin
        _zz_shift_q_7 = shift_q_map_16;
      end
      6'b010001 : begin
        _zz_shift_q_7 = shift_q_map_17;
      end
      6'b010010 : begin
        _zz_shift_q_7 = shift_q_map_18;
      end
      6'b010011 : begin
        _zz_shift_q_7 = shift_q_map_19;
      end
      6'b010100 : begin
        _zz_shift_q_7 = shift_q_map_20;
      end
      6'b010101 : begin
        _zz_shift_q_7 = shift_q_map_21;
      end
      6'b010110 : begin
        _zz_shift_q_7 = shift_q_map_22;
      end
      6'b010111 : begin
        _zz_shift_q_7 = shift_q_map_23;
      end
      6'b011000 : begin
        _zz_shift_q_7 = shift_q_map_24;
      end
      6'b011001 : begin
        _zz_shift_q_7 = shift_q_map_25;
      end
      6'b011010 : begin
        _zz_shift_q_7 = shift_q_map_26;
      end
      6'b011011 : begin
        _zz_shift_q_7 = shift_q_map_27;
      end
      6'b011100 : begin
        _zz_shift_q_7 = shift_q_map_28;
      end
      6'b011101 : begin
        _zz_shift_q_7 = shift_q_map_29;
      end
      6'b011110 : begin
        _zz_shift_q_7 = shift_q_map_30;
      end
      6'b011111 : begin
        _zz_shift_q_7 = shift_q_map_31;
      end
      6'b100000 : begin
        _zz_shift_q_7 = shift_q_map_32;
      end
      6'b100001 : begin
        _zz_shift_q_7 = shift_q_map_33;
      end
      6'b100010 : begin
        _zz_shift_q_7 = shift_q_map_34;
      end
      6'b100011 : begin
        _zz_shift_q_7 = shift_q_map_35;
      end
      6'b100100 : begin
        _zz_shift_q_7 = shift_q_map_36;
      end
      6'b100101 : begin
        _zz_shift_q_7 = shift_q_map_37;
      end
      6'b100110 : begin
        _zz_shift_q_7 = shift_q_map_38;
      end
      default : begin
        _zz_shift_q_7 = shift_q_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_0_3)
      6'b000000 : begin
        _zz_shift_i_0_2 = shift_i_map_0;
      end
      6'b000001 : begin
        _zz_shift_i_0_2 = shift_i_map_1;
      end
      6'b000010 : begin
        _zz_shift_i_0_2 = shift_i_map_2;
      end
      6'b000011 : begin
        _zz_shift_i_0_2 = shift_i_map_3;
      end
      6'b000100 : begin
        _zz_shift_i_0_2 = shift_i_map_4;
      end
      6'b000101 : begin
        _zz_shift_i_0_2 = shift_i_map_5;
      end
      6'b000110 : begin
        _zz_shift_i_0_2 = shift_i_map_6;
      end
      6'b000111 : begin
        _zz_shift_i_0_2 = shift_i_map_7;
      end
      6'b001000 : begin
        _zz_shift_i_0_2 = shift_i_map_8;
      end
      6'b001001 : begin
        _zz_shift_i_0_2 = shift_i_map_9;
      end
      6'b001010 : begin
        _zz_shift_i_0_2 = shift_i_map_10;
      end
      6'b001011 : begin
        _zz_shift_i_0_2 = shift_i_map_11;
      end
      6'b001100 : begin
        _zz_shift_i_0_2 = shift_i_map_12;
      end
      6'b001101 : begin
        _zz_shift_i_0_2 = shift_i_map_13;
      end
      6'b001110 : begin
        _zz_shift_i_0_2 = shift_i_map_14;
      end
      6'b001111 : begin
        _zz_shift_i_0_2 = shift_i_map_15;
      end
      6'b010000 : begin
        _zz_shift_i_0_2 = shift_i_map_16;
      end
      6'b010001 : begin
        _zz_shift_i_0_2 = shift_i_map_17;
      end
      6'b010010 : begin
        _zz_shift_i_0_2 = shift_i_map_18;
      end
      6'b010011 : begin
        _zz_shift_i_0_2 = shift_i_map_19;
      end
      6'b010100 : begin
        _zz_shift_i_0_2 = shift_i_map_20;
      end
      6'b010101 : begin
        _zz_shift_i_0_2 = shift_i_map_21;
      end
      6'b010110 : begin
        _zz_shift_i_0_2 = shift_i_map_22;
      end
      6'b010111 : begin
        _zz_shift_i_0_2 = shift_i_map_23;
      end
      6'b011000 : begin
        _zz_shift_i_0_2 = shift_i_map_24;
      end
      6'b011001 : begin
        _zz_shift_i_0_2 = shift_i_map_25;
      end
      6'b011010 : begin
        _zz_shift_i_0_2 = shift_i_map_26;
      end
      6'b011011 : begin
        _zz_shift_i_0_2 = shift_i_map_27;
      end
      6'b011100 : begin
        _zz_shift_i_0_2 = shift_i_map_28;
      end
      6'b011101 : begin
        _zz_shift_i_0_2 = shift_i_map_29;
      end
      6'b011110 : begin
        _zz_shift_i_0_2 = shift_i_map_30;
      end
      6'b011111 : begin
        _zz_shift_i_0_2 = shift_i_map_31;
      end
      6'b100000 : begin
        _zz_shift_i_0_2 = shift_i_map_32;
      end
      6'b100001 : begin
        _zz_shift_i_0_2 = shift_i_map_33;
      end
      6'b100010 : begin
        _zz_shift_i_0_2 = shift_i_map_34;
      end
      6'b100011 : begin
        _zz_shift_i_0_2 = shift_i_map_35;
      end
      6'b100100 : begin
        _zz_shift_i_0_2 = shift_i_map_36;
      end
      6'b100101 : begin
        _zz_shift_i_0_2 = shift_i_map_37;
      end
      6'b100110 : begin
        _zz_shift_i_0_2 = shift_i_map_38;
      end
      default : begin
        _zz_shift_i_0_2 = shift_i_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_0_3)
      6'b000000 : begin
        _zz_shift_q_0_2 = shift_q_map_0;
      end
      6'b000001 : begin
        _zz_shift_q_0_2 = shift_q_map_1;
      end
      6'b000010 : begin
        _zz_shift_q_0_2 = shift_q_map_2;
      end
      6'b000011 : begin
        _zz_shift_q_0_2 = shift_q_map_3;
      end
      6'b000100 : begin
        _zz_shift_q_0_2 = shift_q_map_4;
      end
      6'b000101 : begin
        _zz_shift_q_0_2 = shift_q_map_5;
      end
      6'b000110 : begin
        _zz_shift_q_0_2 = shift_q_map_6;
      end
      6'b000111 : begin
        _zz_shift_q_0_2 = shift_q_map_7;
      end
      6'b001000 : begin
        _zz_shift_q_0_2 = shift_q_map_8;
      end
      6'b001001 : begin
        _zz_shift_q_0_2 = shift_q_map_9;
      end
      6'b001010 : begin
        _zz_shift_q_0_2 = shift_q_map_10;
      end
      6'b001011 : begin
        _zz_shift_q_0_2 = shift_q_map_11;
      end
      6'b001100 : begin
        _zz_shift_q_0_2 = shift_q_map_12;
      end
      6'b001101 : begin
        _zz_shift_q_0_2 = shift_q_map_13;
      end
      6'b001110 : begin
        _zz_shift_q_0_2 = shift_q_map_14;
      end
      6'b001111 : begin
        _zz_shift_q_0_2 = shift_q_map_15;
      end
      6'b010000 : begin
        _zz_shift_q_0_2 = shift_q_map_16;
      end
      6'b010001 : begin
        _zz_shift_q_0_2 = shift_q_map_17;
      end
      6'b010010 : begin
        _zz_shift_q_0_2 = shift_q_map_18;
      end
      6'b010011 : begin
        _zz_shift_q_0_2 = shift_q_map_19;
      end
      6'b010100 : begin
        _zz_shift_q_0_2 = shift_q_map_20;
      end
      6'b010101 : begin
        _zz_shift_q_0_2 = shift_q_map_21;
      end
      6'b010110 : begin
        _zz_shift_q_0_2 = shift_q_map_22;
      end
      6'b010111 : begin
        _zz_shift_q_0_2 = shift_q_map_23;
      end
      6'b011000 : begin
        _zz_shift_q_0_2 = shift_q_map_24;
      end
      6'b011001 : begin
        _zz_shift_q_0_2 = shift_q_map_25;
      end
      6'b011010 : begin
        _zz_shift_q_0_2 = shift_q_map_26;
      end
      6'b011011 : begin
        _zz_shift_q_0_2 = shift_q_map_27;
      end
      6'b011100 : begin
        _zz_shift_q_0_2 = shift_q_map_28;
      end
      6'b011101 : begin
        _zz_shift_q_0_2 = shift_q_map_29;
      end
      6'b011110 : begin
        _zz_shift_q_0_2 = shift_q_map_30;
      end
      6'b011111 : begin
        _zz_shift_q_0_2 = shift_q_map_31;
      end
      6'b100000 : begin
        _zz_shift_q_0_2 = shift_q_map_32;
      end
      6'b100001 : begin
        _zz_shift_q_0_2 = shift_q_map_33;
      end
      6'b100010 : begin
        _zz_shift_q_0_2 = shift_q_map_34;
      end
      6'b100011 : begin
        _zz_shift_q_0_2 = shift_q_map_35;
      end
      6'b100100 : begin
        _zz_shift_q_0_2 = shift_q_map_36;
      end
      6'b100101 : begin
        _zz_shift_q_0_2 = shift_q_map_37;
      end
      6'b100110 : begin
        _zz_shift_q_0_2 = shift_q_map_38;
      end
      default : begin
        _zz_shift_q_0_2 = shift_q_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_1_3)
      6'b000000 : begin
        _zz_shift_i_1_2 = shift_i_map_0;
      end
      6'b000001 : begin
        _zz_shift_i_1_2 = shift_i_map_1;
      end
      6'b000010 : begin
        _zz_shift_i_1_2 = shift_i_map_2;
      end
      6'b000011 : begin
        _zz_shift_i_1_2 = shift_i_map_3;
      end
      6'b000100 : begin
        _zz_shift_i_1_2 = shift_i_map_4;
      end
      6'b000101 : begin
        _zz_shift_i_1_2 = shift_i_map_5;
      end
      6'b000110 : begin
        _zz_shift_i_1_2 = shift_i_map_6;
      end
      6'b000111 : begin
        _zz_shift_i_1_2 = shift_i_map_7;
      end
      6'b001000 : begin
        _zz_shift_i_1_2 = shift_i_map_8;
      end
      6'b001001 : begin
        _zz_shift_i_1_2 = shift_i_map_9;
      end
      6'b001010 : begin
        _zz_shift_i_1_2 = shift_i_map_10;
      end
      6'b001011 : begin
        _zz_shift_i_1_2 = shift_i_map_11;
      end
      6'b001100 : begin
        _zz_shift_i_1_2 = shift_i_map_12;
      end
      6'b001101 : begin
        _zz_shift_i_1_2 = shift_i_map_13;
      end
      6'b001110 : begin
        _zz_shift_i_1_2 = shift_i_map_14;
      end
      6'b001111 : begin
        _zz_shift_i_1_2 = shift_i_map_15;
      end
      6'b010000 : begin
        _zz_shift_i_1_2 = shift_i_map_16;
      end
      6'b010001 : begin
        _zz_shift_i_1_2 = shift_i_map_17;
      end
      6'b010010 : begin
        _zz_shift_i_1_2 = shift_i_map_18;
      end
      6'b010011 : begin
        _zz_shift_i_1_2 = shift_i_map_19;
      end
      6'b010100 : begin
        _zz_shift_i_1_2 = shift_i_map_20;
      end
      6'b010101 : begin
        _zz_shift_i_1_2 = shift_i_map_21;
      end
      6'b010110 : begin
        _zz_shift_i_1_2 = shift_i_map_22;
      end
      6'b010111 : begin
        _zz_shift_i_1_2 = shift_i_map_23;
      end
      6'b011000 : begin
        _zz_shift_i_1_2 = shift_i_map_24;
      end
      6'b011001 : begin
        _zz_shift_i_1_2 = shift_i_map_25;
      end
      6'b011010 : begin
        _zz_shift_i_1_2 = shift_i_map_26;
      end
      6'b011011 : begin
        _zz_shift_i_1_2 = shift_i_map_27;
      end
      6'b011100 : begin
        _zz_shift_i_1_2 = shift_i_map_28;
      end
      6'b011101 : begin
        _zz_shift_i_1_2 = shift_i_map_29;
      end
      6'b011110 : begin
        _zz_shift_i_1_2 = shift_i_map_30;
      end
      6'b011111 : begin
        _zz_shift_i_1_2 = shift_i_map_31;
      end
      6'b100000 : begin
        _zz_shift_i_1_2 = shift_i_map_32;
      end
      6'b100001 : begin
        _zz_shift_i_1_2 = shift_i_map_33;
      end
      6'b100010 : begin
        _zz_shift_i_1_2 = shift_i_map_34;
      end
      6'b100011 : begin
        _zz_shift_i_1_2 = shift_i_map_35;
      end
      6'b100100 : begin
        _zz_shift_i_1_2 = shift_i_map_36;
      end
      6'b100101 : begin
        _zz_shift_i_1_2 = shift_i_map_37;
      end
      6'b100110 : begin
        _zz_shift_i_1_2 = shift_i_map_38;
      end
      default : begin
        _zz_shift_i_1_2 = shift_i_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_1_3)
      6'b000000 : begin
        _zz_shift_q_1_2 = shift_q_map_0;
      end
      6'b000001 : begin
        _zz_shift_q_1_2 = shift_q_map_1;
      end
      6'b000010 : begin
        _zz_shift_q_1_2 = shift_q_map_2;
      end
      6'b000011 : begin
        _zz_shift_q_1_2 = shift_q_map_3;
      end
      6'b000100 : begin
        _zz_shift_q_1_2 = shift_q_map_4;
      end
      6'b000101 : begin
        _zz_shift_q_1_2 = shift_q_map_5;
      end
      6'b000110 : begin
        _zz_shift_q_1_2 = shift_q_map_6;
      end
      6'b000111 : begin
        _zz_shift_q_1_2 = shift_q_map_7;
      end
      6'b001000 : begin
        _zz_shift_q_1_2 = shift_q_map_8;
      end
      6'b001001 : begin
        _zz_shift_q_1_2 = shift_q_map_9;
      end
      6'b001010 : begin
        _zz_shift_q_1_2 = shift_q_map_10;
      end
      6'b001011 : begin
        _zz_shift_q_1_2 = shift_q_map_11;
      end
      6'b001100 : begin
        _zz_shift_q_1_2 = shift_q_map_12;
      end
      6'b001101 : begin
        _zz_shift_q_1_2 = shift_q_map_13;
      end
      6'b001110 : begin
        _zz_shift_q_1_2 = shift_q_map_14;
      end
      6'b001111 : begin
        _zz_shift_q_1_2 = shift_q_map_15;
      end
      6'b010000 : begin
        _zz_shift_q_1_2 = shift_q_map_16;
      end
      6'b010001 : begin
        _zz_shift_q_1_2 = shift_q_map_17;
      end
      6'b010010 : begin
        _zz_shift_q_1_2 = shift_q_map_18;
      end
      6'b010011 : begin
        _zz_shift_q_1_2 = shift_q_map_19;
      end
      6'b010100 : begin
        _zz_shift_q_1_2 = shift_q_map_20;
      end
      6'b010101 : begin
        _zz_shift_q_1_2 = shift_q_map_21;
      end
      6'b010110 : begin
        _zz_shift_q_1_2 = shift_q_map_22;
      end
      6'b010111 : begin
        _zz_shift_q_1_2 = shift_q_map_23;
      end
      6'b011000 : begin
        _zz_shift_q_1_2 = shift_q_map_24;
      end
      6'b011001 : begin
        _zz_shift_q_1_2 = shift_q_map_25;
      end
      6'b011010 : begin
        _zz_shift_q_1_2 = shift_q_map_26;
      end
      6'b011011 : begin
        _zz_shift_q_1_2 = shift_q_map_27;
      end
      6'b011100 : begin
        _zz_shift_q_1_2 = shift_q_map_28;
      end
      6'b011101 : begin
        _zz_shift_q_1_2 = shift_q_map_29;
      end
      6'b011110 : begin
        _zz_shift_q_1_2 = shift_q_map_30;
      end
      6'b011111 : begin
        _zz_shift_q_1_2 = shift_q_map_31;
      end
      6'b100000 : begin
        _zz_shift_q_1_2 = shift_q_map_32;
      end
      6'b100001 : begin
        _zz_shift_q_1_2 = shift_q_map_33;
      end
      6'b100010 : begin
        _zz_shift_q_1_2 = shift_q_map_34;
      end
      6'b100011 : begin
        _zz_shift_q_1_2 = shift_q_map_35;
      end
      6'b100100 : begin
        _zz_shift_q_1_2 = shift_q_map_36;
      end
      6'b100101 : begin
        _zz_shift_q_1_2 = shift_q_map_37;
      end
      6'b100110 : begin
        _zz_shift_q_1_2 = shift_q_map_38;
      end
      default : begin
        _zz_shift_q_1_2 = shift_q_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_2_3)
      6'b000000 : begin
        _zz_shift_i_2_2 = shift_i_map_0;
      end
      6'b000001 : begin
        _zz_shift_i_2_2 = shift_i_map_1;
      end
      6'b000010 : begin
        _zz_shift_i_2_2 = shift_i_map_2;
      end
      6'b000011 : begin
        _zz_shift_i_2_2 = shift_i_map_3;
      end
      6'b000100 : begin
        _zz_shift_i_2_2 = shift_i_map_4;
      end
      6'b000101 : begin
        _zz_shift_i_2_2 = shift_i_map_5;
      end
      6'b000110 : begin
        _zz_shift_i_2_2 = shift_i_map_6;
      end
      6'b000111 : begin
        _zz_shift_i_2_2 = shift_i_map_7;
      end
      6'b001000 : begin
        _zz_shift_i_2_2 = shift_i_map_8;
      end
      6'b001001 : begin
        _zz_shift_i_2_2 = shift_i_map_9;
      end
      6'b001010 : begin
        _zz_shift_i_2_2 = shift_i_map_10;
      end
      6'b001011 : begin
        _zz_shift_i_2_2 = shift_i_map_11;
      end
      6'b001100 : begin
        _zz_shift_i_2_2 = shift_i_map_12;
      end
      6'b001101 : begin
        _zz_shift_i_2_2 = shift_i_map_13;
      end
      6'b001110 : begin
        _zz_shift_i_2_2 = shift_i_map_14;
      end
      6'b001111 : begin
        _zz_shift_i_2_2 = shift_i_map_15;
      end
      6'b010000 : begin
        _zz_shift_i_2_2 = shift_i_map_16;
      end
      6'b010001 : begin
        _zz_shift_i_2_2 = shift_i_map_17;
      end
      6'b010010 : begin
        _zz_shift_i_2_2 = shift_i_map_18;
      end
      6'b010011 : begin
        _zz_shift_i_2_2 = shift_i_map_19;
      end
      6'b010100 : begin
        _zz_shift_i_2_2 = shift_i_map_20;
      end
      6'b010101 : begin
        _zz_shift_i_2_2 = shift_i_map_21;
      end
      6'b010110 : begin
        _zz_shift_i_2_2 = shift_i_map_22;
      end
      6'b010111 : begin
        _zz_shift_i_2_2 = shift_i_map_23;
      end
      6'b011000 : begin
        _zz_shift_i_2_2 = shift_i_map_24;
      end
      6'b011001 : begin
        _zz_shift_i_2_2 = shift_i_map_25;
      end
      6'b011010 : begin
        _zz_shift_i_2_2 = shift_i_map_26;
      end
      6'b011011 : begin
        _zz_shift_i_2_2 = shift_i_map_27;
      end
      6'b011100 : begin
        _zz_shift_i_2_2 = shift_i_map_28;
      end
      6'b011101 : begin
        _zz_shift_i_2_2 = shift_i_map_29;
      end
      6'b011110 : begin
        _zz_shift_i_2_2 = shift_i_map_30;
      end
      6'b011111 : begin
        _zz_shift_i_2_2 = shift_i_map_31;
      end
      6'b100000 : begin
        _zz_shift_i_2_2 = shift_i_map_32;
      end
      6'b100001 : begin
        _zz_shift_i_2_2 = shift_i_map_33;
      end
      6'b100010 : begin
        _zz_shift_i_2_2 = shift_i_map_34;
      end
      6'b100011 : begin
        _zz_shift_i_2_2 = shift_i_map_35;
      end
      6'b100100 : begin
        _zz_shift_i_2_2 = shift_i_map_36;
      end
      6'b100101 : begin
        _zz_shift_i_2_2 = shift_i_map_37;
      end
      6'b100110 : begin
        _zz_shift_i_2_2 = shift_i_map_38;
      end
      default : begin
        _zz_shift_i_2_2 = shift_i_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_2_3)
      6'b000000 : begin
        _zz_shift_q_2_2 = shift_q_map_0;
      end
      6'b000001 : begin
        _zz_shift_q_2_2 = shift_q_map_1;
      end
      6'b000010 : begin
        _zz_shift_q_2_2 = shift_q_map_2;
      end
      6'b000011 : begin
        _zz_shift_q_2_2 = shift_q_map_3;
      end
      6'b000100 : begin
        _zz_shift_q_2_2 = shift_q_map_4;
      end
      6'b000101 : begin
        _zz_shift_q_2_2 = shift_q_map_5;
      end
      6'b000110 : begin
        _zz_shift_q_2_2 = shift_q_map_6;
      end
      6'b000111 : begin
        _zz_shift_q_2_2 = shift_q_map_7;
      end
      6'b001000 : begin
        _zz_shift_q_2_2 = shift_q_map_8;
      end
      6'b001001 : begin
        _zz_shift_q_2_2 = shift_q_map_9;
      end
      6'b001010 : begin
        _zz_shift_q_2_2 = shift_q_map_10;
      end
      6'b001011 : begin
        _zz_shift_q_2_2 = shift_q_map_11;
      end
      6'b001100 : begin
        _zz_shift_q_2_2 = shift_q_map_12;
      end
      6'b001101 : begin
        _zz_shift_q_2_2 = shift_q_map_13;
      end
      6'b001110 : begin
        _zz_shift_q_2_2 = shift_q_map_14;
      end
      6'b001111 : begin
        _zz_shift_q_2_2 = shift_q_map_15;
      end
      6'b010000 : begin
        _zz_shift_q_2_2 = shift_q_map_16;
      end
      6'b010001 : begin
        _zz_shift_q_2_2 = shift_q_map_17;
      end
      6'b010010 : begin
        _zz_shift_q_2_2 = shift_q_map_18;
      end
      6'b010011 : begin
        _zz_shift_q_2_2 = shift_q_map_19;
      end
      6'b010100 : begin
        _zz_shift_q_2_2 = shift_q_map_20;
      end
      6'b010101 : begin
        _zz_shift_q_2_2 = shift_q_map_21;
      end
      6'b010110 : begin
        _zz_shift_q_2_2 = shift_q_map_22;
      end
      6'b010111 : begin
        _zz_shift_q_2_2 = shift_q_map_23;
      end
      6'b011000 : begin
        _zz_shift_q_2_2 = shift_q_map_24;
      end
      6'b011001 : begin
        _zz_shift_q_2_2 = shift_q_map_25;
      end
      6'b011010 : begin
        _zz_shift_q_2_2 = shift_q_map_26;
      end
      6'b011011 : begin
        _zz_shift_q_2_2 = shift_q_map_27;
      end
      6'b011100 : begin
        _zz_shift_q_2_2 = shift_q_map_28;
      end
      6'b011101 : begin
        _zz_shift_q_2_2 = shift_q_map_29;
      end
      6'b011110 : begin
        _zz_shift_q_2_2 = shift_q_map_30;
      end
      6'b011111 : begin
        _zz_shift_q_2_2 = shift_q_map_31;
      end
      6'b100000 : begin
        _zz_shift_q_2_2 = shift_q_map_32;
      end
      6'b100001 : begin
        _zz_shift_q_2_2 = shift_q_map_33;
      end
      6'b100010 : begin
        _zz_shift_q_2_2 = shift_q_map_34;
      end
      6'b100011 : begin
        _zz_shift_q_2_2 = shift_q_map_35;
      end
      6'b100100 : begin
        _zz_shift_q_2_2 = shift_q_map_36;
      end
      6'b100101 : begin
        _zz_shift_q_2_2 = shift_q_map_37;
      end
      6'b100110 : begin
        _zz_shift_q_2_2 = shift_q_map_38;
      end
      default : begin
        _zz_shift_q_2_2 = shift_q_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_3_3)
      6'b000000 : begin
        _zz_shift_i_3_2 = shift_i_map_0;
      end
      6'b000001 : begin
        _zz_shift_i_3_2 = shift_i_map_1;
      end
      6'b000010 : begin
        _zz_shift_i_3_2 = shift_i_map_2;
      end
      6'b000011 : begin
        _zz_shift_i_3_2 = shift_i_map_3;
      end
      6'b000100 : begin
        _zz_shift_i_3_2 = shift_i_map_4;
      end
      6'b000101 : begin
        _zz_shift_i_3_2 = shift_i_map_5;
      end
      6'b000110 : begin
        _zz_shift_i_3_2 = shift_i_map_6;
      end
      6'b000111 : begin
        _zz_shift_i_3_2 = shift_i_map_7;
      end
      6'b001000 : begin
        _zz_shift_i_3_2 = shift_i_map_8;
      end
      6'b001001 : begin
        _zz_shift_i_3_2 = shift_i_map_9;
      end
      6'b001010 : begin
        _zz_shift_i_3_2 = shift_i_map_10;
      end
      6'b001011 : begin
        _zz_shift_i_3_2 = shift_i_map_11;
      end
      6'b001100 : begin
        _zz_shift_i_3_2 = shift_i_map_12;
      end
      6'b001101 : begin
        _zz_shift_i_3_2 = shift_i_map_13;
      end
      6'b001110 : begin
        _zz_shift_i_3_2 = shift_i_map_14;
      end
      6'b001111 : begin
        _zz_shift_i_3_2 = shift_i_map_15;
      end
      6'b010000 : begin
        _zz_shift_i_3_2 = shift_i_map_16;
      end
      6'b010001 : begin
        _zz_shift_i_3_2 = shift_i_map_17;
      end
      6'b010010 : begin
        _zz_shift_i_3_2 = shift_i_map_18;
      end
      6'b010011 : begin
        _zz_shift_i_3_2 = shift_i_map_19;
      end
      6'b010100 : begin
        _zz_shift_i_3_2 = shift_i_map_20;
      end
      6'b010101 : begin
        _zz_shift_i_3_2 = shift_i_map_21;
      end
      6'b010110 : begin
        _zz_shift_i_3_2 = shift_i_map_22;
      end
      6'b010111 : begin
        _zz_shift_i_3_2 = shift_i_map_23;
      end
      6'b011000 : begin
        _zz_shift_i_3_2 = shift_i_map_24;
      end
      6'b011001 : begin
        _zz_shift_i_3_2 = shift_i_map_25;
      end
      6'b011010 : begin
        _zz_shift_i_3_2 = shift_i_map_26;
      end
      6'b011011 : begin
        _zz_shift_i_3_2 = shift_i_map_27;
      end
      6'b011100 : begin
        _zz_shift_i_3_2 = shift_i_map_28;
      end
      6'b011101 : begin
        _zz_shift_i_3_2 = shift_i_map_29;
      end
      6'b011110 : begin
        _zz_shift_i_3_2 = shift_i_map_30;
      end
      6'b011111 : begin
        _zz_shift_i_3_2 = shift_i_map_31;
      end
      6'b100000 : begin
        _zz_shift_i_3_2 = shift_i_map_32;
      end
      6'b100001 : begin
        _zz_shift_i_3_2 = shift_i_map_33;
      end
      6'b100010 : begin
        _zz_shift_i_3_2 = shift_i_map_34;
      end
      6'b100011 : begin
        _zz_shift_i_3_2 = shift_i_map_35;
      end
      6'b100100 : begin
        _zz_shift_i_3_2 = shift_i_map_36;
      end
      6'b100101 : begin
        _zz_shift_i_3_2 = shift_i_map_37;
      end
      6'b100110 : begin
        _zz_shift_i_3_2 = shift_i_map_38;
      end
      default : begin
        _zz_shift_i_3_2 = shift_i_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_3_3)
      6'b000000 : begin
        _zz_shift_q_3_2 = shift_q_map_0;
      end
      6'b000001 : begin
        _zz_shift_q_3_2 = shift_q_map_1;
      end
      6'b000010 : begin
        _zz_shift_q_3_2 = shift_q_map_2;
      end
      6'b000011 : begin
        _zz_shift_q_3_2 = shift_q_map_3;
      end
      6'b000100 : begin
        _zz_shift_q_3_2 = shift_q_map_4;
      end
      6'b000101 : begin
        _zz_shift_q_3_2 = shift_q_map_5;
      end
      6'b000110 : begin
        _zz_shift_q_3_2 = shift_q_map_6;
      end
      6'b000111 : begin
        _zz_shift_q_3_2 = shift_q_map_7;
      end
      6'b001000 : begin
        _zz_shift_q_3_2 = shift_q_map_8;
      end
      6'b001001 : begin
        _zz_shift_q_3_2 = shift_q_map_9;
      end
      6'b001010 : begin
        _zz_shift_q_3_2 = shift_q_map_10;
      end
      6'b001011 : begin
        _zz_shift_q_3_2 = shift_q_map_11;
      end
      6'b001100 : begin
        _zz_shift_q_3_2 = shift_q_map_12;
      end
      6'b001101 : begin
        _zz_shift_q_3_2 = shift_q_map_13;
      end
      6'b001110 : begin
        _zz_shift_q_3_2 = shift_q_map_14;
      end
      6'b001111 : begin
        _zz_shift_q_3_2 = shift_q_map_15;
      end
      6'b010000 : begin
        _zz_shift_q_3_2 = shift_q_map_16;
      end
      6'b010001 : begin
        _zz_shift_q_3_2 = shift_q_map_17;
      end
      6'b010010 : begin
        _zz_shift_q_3_2 = shift_q_map_18;
      end
      6'b010011 : begin
        _zz_shift_q_3_2 = shift_q_map_19;
      end
      6'b010100 : begin
        _zz_shift_q_3_2 = shift_q_map_20;
      end
      6'b010101 : begin
        _zz_shift_q_3_2 = shift_q_map_21;
      end
      6'b010110 : begin
        _zz_shift_q_3_2 = shift_q_map_22;
      end
      6'b010111 : begin
        _zz_shift_q_3_2 = shift_q_map_23;
      end
      6'b011000 : begin
        _zz_shift_q_3_2 = shift_q_map_24;
      end
      6'b011001 : begin
        _zz_shift_q_3_2 = shift_q_map_25;
      end
      6'b011010 : begin
        _zz_shift_q_3_2 = shift_q_map_26;
      end
      6'b011011 : begin
        _zz_shift_q_3_2 = shift_q_map_27;
      end
      6'b011100 : begin
        _zz_shift_q_3_2 = shift_q_map_28;
      end
      6'b011101 : begin
        _zz_shift_q_3_2 = shift_q_map_29;
      end
      6'b011110 : begin
        _zz_shift_q_3_2 = shift_q_map_30;
      end
      6'b011111 : begin
        _zz_shift_q_3_2 = shift_q_map_31;
      end
      6'b100000 : begin
        _zz_shift_q_3_2 = shift_q_map_32;
      end
      6'b100001 : begin
        _zz_shift_q_3_2 = shift_q_map_33;
      end
      6'b100010 : begin
        _zz_shift_q_3_2 = shift_q_map_34;
      end
      6'b100011 : begin
        _zz_shift_q_3_2 = shift_q_map_35;
      end
      6'b100100 : begin
        _zz_shift_q_3_2 = shift_q_map_36;
      end
      6'b100101 : begin
        _zz_shift_q_3_2 = shift_q_map_37;
      end
      6'b100110 : begin
        _zz_shift_q_3_2 = shift_q_map_38;
      end
      default : begin
        _zz_shift_q_3_2 = shift_q_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_4_3)
      6'b000000 : begin
        _zz_shift_i_4_2 = shift_i_map_0;
      end
      6'b000001 : begin
        _zz_shift_i_4_2 = shift_i_map_1;
      end
      6'b000010 : begin
        _zz_shift_i_4_2 = shift_i_map_2;
      end
      6'b000011 : begin
        _zz_shift_i_4_2 = shift_i_map_3;
      end
      6'b000100 : begin
        _zz_shift_i_4_2 = shift_i_map_4;
      end
      6'b000101 : begin
        _zz_shift_i_4_2 = shift_i_map_5;
      end
      6'b000110 : begin
        _zz_shift_i_4_2 = shift_i_map_6;
      end
      6'b000111 : begin
        _zz_shift_i_4_2 = shift_i_map_7;
      end
      6'b001000 : begin
        _zz_shift_i_4_2 = shift_i_map_8;
      end
      6'b001001 : begin
        _zz_shift_i_4_2 = shift_i_map_9;
      end
      6'b001010 : begin
        _zz_shift_i_4_2 = shift_i_map_10;
      end
      6'b001011 : begin
        _zz_shift_i_4_2 = shift_i_map_11;
      end
      6'b001100 : begin
        _zz_shift_i_4_2 = shift_i_map_12;
      end
      6'b001101 : begin
        _zz_shift_i_4_2 = shift_i_map_13;
      end
      6'b001110 : begin
        _zz_shift_i_4_2 = shift_i_map_14;
      end
      6'b001111 : begin
        _zz_shift_i_4_2 = shift_i_map_15;
      end
      6'b010000 : begin
        _zz_shift_i_4_2 = shift_i_map_16;
      end
      6'b010001 : begin
        _zz_shift_i_4_2 = shift_i_map_17;
      end
      6'b010010 : begin
        _zz_shift_i_4_2 = shift_i_map_18;
      end
      6'b010011 : begin
        _zz_shift_i_4_2 = shift_i_map_19;
      end
      6'b010100 : begin
        _zz_shift_i_4_2 = shift_i_map_20;
      end
      6'b010101 : begin
        _zz_shift_i_4_2 = shift_i_map_21;
      end
      6'b010110 : begin
        _zz_shift_i_4_2 = shift_i_map_22;
      end
      6'b010111 : begin
        _zz_shift_i_4_2 = shift_i_map_23;
      end
      6'b011000 : begin
        _zz_shift_i_4_2 = shift_i_map_24;
      end
      6'b011001 : begin
        _zz_shift_i_4_2 = shift_i_map_25;
      end
      6'b011010 : begin
        _zz_shift_i_4_2 = shift_i_map_26;
      end
      6'b011011 : begin
        _zz_shift_i_4_2 = shift_i_map_27;
      end
      6'b011100 : begin
        _zz_shift_i_4_2 = shift_i_map_28;
      end
      6'b011101 : begin
        _zz_shift_i_4_2 = shift_i_map_29;
      end
      6'b011110 : begin
        _zz_shift_i_4_2 = shift_i_map_30;
      end
      6'b011111 : begin
        _zz_shift_i_4_2 = shift_i_map_31;
      end
      6'b100000 : begin
        _zz_shift_i_4_2 = shift_i_map_32;
      end
      6'b100001 : begin
        _zz_shift_i_4_2 = shift_i_map_33;
      end
      6'b100010 : begin
        _zz_shift_i_4_2 = shift_i_map_34;
      end
      6'b100011 : begin
        _zz_shift_i_4_2 = shift_i_map_35;
      end
      6'b100100 : begin
        _zz_shift_i_4_2 = shift_i_map_36;
      end
      6'b100101 : begin
        _zz_shift_i_4_2 = shift_i_map_37;
      end
      6'b100110 : begin
        _zz_shift_i_4_2 = shift_i_map_38;
      end
      default : begin
        _zz_shift_i_4_2 = shift_i_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_4_3)
      6'b000000 : begin
        _zz_shift_q_4_2 = shift_q_map_0;
      end
      6'b000001 : begin
        _zz_shift_q_4_2 = shift_q_map_1;
      end
      6'b000010 : begin
        _zz_shift_q_4_2 = shift_q_map_2;
      end
      6'b000011 : begin
        _zz_shift_q_4_2 = shift_q_map_3;
      end
      6'b000100 : begin
        _zz_shift_q_4_2 = shift_q_map_4;
      end
      6'b000101 : begin
        _zz_shift_q_4_2 = shift_q_map_5;
      end
      6'b000110 : begin
        _zz_shift_q_4_2 = shift_q_map_6;
      end
      6'b000111 : begin
        _zz_shift_q_4_2 = shift_q_map_7;
      end
      6'b001000 : begin
        _zz_shift_q_4_2 = shift_q_map_8;
      end
      6'b001001 : begin
        _zz_shift_q_4_2 = shift_q_map_9;
      end
      6'b001010 : begin
        _zz_shift_q_4_2 = shift_q_map_10;
      end
      6'b001011 : begin
        _zz_shift_q_4_2 = shift_q_map_11;
      end
      6'b001100 : begin
        _zz_shift_q_4_2 = shift_q_map_12;
      end
      6'b001101 : begin
        _zz_shift_q_4_2 = shift_q_map_13;
      end
      6'b001110 : begin
        _zz_shift_q_4_2 = shift_q_map_14;
      end
      6'b001111 : begin
        _zz_shift_q_4_2 = shift_q_map_15;
      end
      6'b010000 : begin
        _zz_shift_q_4_2 = shift_q_map_16;
      end
      6'b010001 : begin
        _zz_shift_q_4_2 = shift_q_map_17;
      end
      6'b010010 : begin
        _zz_shift_q_4_2 = shift_q_map_18;
      end
      6'b010011 : begin
        _zz_shift_q_4_2 = shift_q_map_19;
      end
      6'b010100 : begin
        _zz_shift_q_4_2 = shift_q_map_20;
      end
      6'b010101 : begin
        _zz_shift_q_4_2 = shift_q_map_21;
      end
      6'b010110 : begin
        _zz_shift_q_4_2 = shift_q_map_22;
      end
      6'b010111 : begin
        _zz_shift_q_4_2 = shift_q_map_23;
      end
      6'b011000 : begin
        _zz_shift_q_4_2 = shift_q_map_24;
      end
      6'b011001 : begin
        _zz_shift_q_4_2 = shift_q_map_25;
      end
      6'b011010 : begin
        _zz_shift_q_4_2 = shift_q_map_26;
      end
      6'b011011 : begin
        _zz_shift_q_4_2 = shift_q_map_27;
      end
      6'b011100 : begin
        _zz_shift_q_4_2 = shift_q_map_28;
      end
      6'b011101 : begin
        _zz_shift_q_4_2 = shift_q_map_29;
      end
      6'b011110 : begin
        _zz_shift_q_4_2 = shift_q_map_30;
      end
      6'b011111 : begin
        _zz_shift_q_4_2 = shift_q_map_31;
      end
      6'b100000 : begin
        _zz_shift_q_4_2 = shift_q_map_32;
      end
      6'b100001 : begin
        _zz_shift_q_4_2 = shift_q_map_33;
      end
      6'b100010 : begin
        _zz_shift_q_4_2 = shift_q_map_34;
      end
      6'b100011 : begin
        _zz_shift_q_4_2 = shift_q_map_35;
      end
      6'b100100 : begin
        _zz_shift_q_4_2 = shift_q_map_36;
      end
      6'b100101 : begin
        _zz_shift_q_4_2 = shift_q_map_37;
      end
      6'b100110 : begin
        _zz_shift_q_4_2 = shift_q_map_38;
      end
      default : begin
        _zz_shift_q_4_2 = shift_q_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_5_3)
      6'b000000 : begin
        _zz_shift_i_5_2 = shift_i_map_0;
      end
      6'b000001 : begin
        _zz_shift_i_5_2 = shift_i_map_1;
      end
      6'b000010 : begin
        _zz_shift_i_5_2 = shift_i_map_2;
      end
      6'b000011 : begin
        _zz_shift_i_5_2 = shift_i_map_3;
      end
      6'b000100 : begin
        _zz_shift_i_5_2 = shift_i_map_4;
      end
      6'b000101 : begin
        _zz_shift_i_5_2 = shift_i_map_5;
      end
      6'b000110 : begin
        _zz_shift_i_5_2 = shift_i_map_6;
      end
      6'b000111 : begin
        _zz_shift_i_5_2 = shift_i_map_7;
      end
      6'b001000 : begin
        _zz_shift_i_5_2 = shift_i_map_8;
      end
      6'b001001 : begin
        _zz_shift_i_5_2 = shift_i_map_9;
      end
      6'b001010 : begin
        _zz_shift_i_5_2 = shift_i_map_10;
      end
      6'b001011 : begin
        _zz_shift_i_5_2 = shift_i_map_11;
      end
      6'b001100 : begin
        _zz_shift_i_5_2 = shift_i_map_12;
      end
      6'b001101 : begin
        _zz_shift_i_5_2 = shift_i_map_13;
      end
      6'b001110 : begin
        _zz_shift_i_5_2 = shift_i_map_14;
      end
      6'b001111 : begin
        _zz_shift_i_5_2 = shift_i_map_15;
      end
      6'b010000 : begin
        _zz_shift_i_5_2 = shift_i_map_16;
      end
      6'b010001 : begin
        _zz_shift_i_5_2 = shift_i_map_17;
      end
      6'b010010 : begin
        _zz_shift_i_5_2 = shift_i_map_18;
      end
      6'b010011 : begin
        _zz_shift_i_5_2 = shift_i_map_19;
      end
      6'b010100 : begin
        _zz_shift_i_5_2 = shift_i_map_20;
      end
      6'b010101 : begin
        _zz_shift_i_5_2 = shift_i_map_21;
      end
      6'b010110 : begin
        _zz_shift_i_5_2 = shift_i_map_22;
      end
      6'b010111 : begin
        _zz_shift_i_5_2 = shift_i_map_23;
      end
      6'b011000 : begin
        _zz_shift_i_5_2 = shift_i_map_24;
      end
      6'b011001 : begin
        _zz_shift_i_5_2 = shift_i_map_25;
      end
      6'b011010 : begin
        _zz_shift_i_5_2 = shift_i_map_26;
      end
      6'b011011 : begin
        _zz_shift_i_5_2 = shift_i_map_27;
      end
      6'b011100 : begin
        _zz_shift_i_5_2 = shift_i_map_28;
      end
      6'b011101 : begin
        _zz_shift_i_5_2 = shift_i_map_29;
      end
      6'b011110 : begin
        _zz_shift_i_5_2 = shift_i_map_30;
      end
      6'b011111 : begin
        _zz_shift_i_5_2 = shift_i_map_31;
      end
      6'b100000 : begin
        _zz_shift_i_5_2 = shift_i_map_32;
      end
      6'b100001 : begin
        _zz_shift_i_5_2 = shift_i_map_33;
      end
      6'b100010 : begin
        _zz_shift_i_5_2 = shift_i_map_34;
      end
      6'b100011 : begin
        _zz_shift_i_5_2 = shift_i_map_35;
      end
      6'b100100 : begin
        _zz_shift_i_5_2 = shift_i_map_36;
      end
      6'b100101 : begin
        _zz_shift_i_5_2 = shift_i_map_37;
      end
      6'b100110 : begin
        _zz_shift_i_5_2 = shift_i_map_38;
      end
      default : begin
        _zz_shift_i_5_2 = shift_i_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_5_3)
      6'b000000 : begin
        _zz_shift_q_5_2 = shift_q_map_0;
      end
      6'b000001 : begin
        _zz_shift_q_5_2 = shift_q_map_1;
      end
      6'b000010 : begin
        _zz_shift_q_5_2 = shift_q_map_2;
      end
      6'b000011 : begin
        _zz_shift_q_5_2 = shift_q_map_3;
      end
      6'b000100 : begin
        _zz_shift_q_5_2 = shift_q_map_4;
      end
      6'b000101 : begin
        _zz_shift_q_5_2 = shift_q_map_5;
      end
      6'b000110 : begin
        _zz_shift_q_5_2 = shift_q_map_6;
      end
      6'b000111 : begin
        _zz_shift_q_5_2 = shift_q_map_7;
      end
      6'b001000 : begin
        _zz_shift_q_5_2 = shift_q_map_8;
      end
      6'b001001 : begin
        _zz_shift_q_5_2 = shift_q_map_9;
      end
      6'b001010 : begin
        _zz_shift_q_5_2 = shift_q_map_10;
      end
      6'b001011 : begin
        _zz_shift_q_5_2 = shift_q_map_11;
      end
      6'b001100 : begin
        _zz_shift_q_5_2 = shift_q_map_12;
      end
      6'b001101 : begin
        _zz_shift_q_5_2 = shift_q_map_13;
      end
      6'b001110 : begin
        _zz_shift_q_5_2 = shift_q_map_14;
      end
      6'b001111 : begin
        _zz_shift_q_5_2 = shift_q_map_15;
      end
      6'b010000 : begin
        _zz_shift_q_5_2 = shift_q_map_16;
      end
      6'b010001 : begin
        _zz_shift_q_5_2 = shift_q_map_17;
      end
      6'b010010 : begin
        _zz_shift_q_5_2 = shift_q_map_18;
      end
      6'b010011 : begin
        _zz_shift_q_5_2 = shift_q_map_19;
      end
      6'b010100 : begin
        _zz_shift_q_5_2 = shift_q_map_20;
      end
      6'b010101 : begin
        _zz_shift_q_5_2 = shift_q_map_21;
      end
      6'b010110 : begin
        _zz_shift_q_5_2 = shift_q_map_22;
      end
      6'b010111 : begin
        _zz_shift_q_5_2 = shift_q_map_23;
      end
      6'b011000 : begin
        _zz_shift_q_5_2 = shift_q_map_24;
      end
      6'b011001 : begin
        _zz_shift_q_5_2 = shift_q_map_25;
      end
      6'b011010 : begin
        _zz_shift_q_5_2 = shift_q_map_26;
      end
      6'b011011 : begin
        _zz_shift_q_5_2 = shift_q_map_27;
      end
      6'b011100 : begin
        _zz_shift_q_5_2 = shift_q_map_28;
      end
      6'b011101 : begin
        _zz_shift_q_5_2 = shift_q_map_29;
      end
      6'b011110 : begin
        _zz_shift_q_5_2 = shift_q_map_30;
      end
      6'b011111 : begin
        _zz_shift_q_5_2 = shift_q_map_31;
      end
      6'b100000 : begin
        _zz_shift_q_5_2 = shift_q_map_32;
      end
      6'b100001 : begin
        _zz_shift_q_5_2 = shift_q_map_33;
      end
      6'b100010 : begin
        _zz_shift_q_5_2 = shift_q_map_34;
      end
      6'b100011 : begin
        _zz_shift_q_5_2 = shift_q_map_35;
      end
      6'b100100 : begin
        _zz_shift_q_5_2 = shift_q_map_36;
      end
      6'b100101 : begin
        _zz_shift_q_5_2 = shift_q_map_37;
      end
      6'b100110 : begin
        _zz_shift_q_5_2 = shift_q_map_38;
      end
      default : begin
        _zz_shift_q_5_2 = shift_q_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_6_3)
      6'b000000 : begin
        _zz_shift_i_6_2 = shift_i_map_0;
      end
      6'b000001 : begin
        _zz_shift_i_6_2 = shift_i_map_1;
      end
      6'b000010 : begin
        _zz_shift_i_6_2 = shift_i_map_2;
      end
      6'b000011 : begin
        _zz_shift_i_6_2 = shift_i_map_3;
      end
      6'b000100 : begin
        _zz_shift_i_6_2 = shift_i_map_4;
      end
      6'b000101 : begin
        _zz_shift_i_6_2 = shift_i_map_5;
      end
      6'b000110 : begin
        _zz_shift_i_6_2 = shift_i_map_6;
      end
      6'b000111 : begin
        _zz_shift_i_6_2 = shift_i_map_7;
      end
      6'b001000 : begin
        _zz_shift_i_6_2 = shift_i_map_8;
      end
      6'b001001 : begin
        _zz_shift_i_6_2 = shift_i_map_9;
      end
      6'b001010 : begin
        _zz_shift_i_6_2 = shift_i_map_10;
      end
      6'b001011 : begin
        _zz_shift_i_6_2 = shift_i_map_11;
      end
      6'b001100 : begin
        _zz_shift_i_6_2 = shift_i_map_12;
      end
      6'b001101 : begin
        _zz_shift_i_6_2 = shift_i_map_13;
      end
      6'b001110 : begin
        _zz_shift_i_6_2 = shift_i_map_14;
      end
      6'b001111 : begin
        _zz_shift_i_6_2 = shift_i_map_15;
      end
      6'b010000 : begin
        _zz_shift_i_6_2 = shift_i_map_16;
      end
      6'b010001 : begin
        _zz_shift_i_6_2 = shift_i_map_17;
      end
      6'b010010 : begin
        _zz_shift_i_6_2 = shift_i_map_18;
      end
      6'b010011 : begin
        _zz_shift_i_6_2 = shift_i_map_19;
      end
      6'b010100 : begin
        _zz_shift_i_6_2 = shift_i_map_20;
      end
      6'b010101 : begin
        _zz_shift_i_6_2 = shift_i_map_21;
      end
      6'b010110 : begin
        _zz_shift_i_6_2 = shift_i_map_22;
      end
      6'b010111 : begin
        _zz_shift_i_6_2 = shift_i_map_23;
      end
      6'b011000 : begin
        _zz_shift_i_6_2 = shift_i_map_24;
      end
      6'b011001 : begin
        _zz_shift_i_6_2 = shift_i_map_25;
      end
      6'b011010 : begin
        _zz_shift_i_6_2 = shift_i_map_26;
      end
      6'b011011 : begin
        _zz_shift_i_6_2 = shift_i_map_27;
      end
      6'b011100 : begin
        _zz_shift_i_6_2 = shift_i_map_28;
      end
      6'b011101 : begin
        _zz_shift_i_6_2 = shift_i_map_29;
      end
      6'b011110 : begin
        _zz_shift_i_6_2 = shift_i_map_30;
      end
      6'b011111 : begin
        _zz_shift_i_6_2 = shift_i_map_31;
      end
      6'b100000 : begin
        _zz_shift_i_6_2 = shift_i_map_32;
      end
      6'b100001 : begin
        _zz_shift_i_6_2 = shift_i_map_33;
      end
      6'b100010 : begin
        _zz_shift_i_6_2 = shift_i_map_34;
      end
      6'b100011 : begin
        _zz_shift_i_6_2 = shift_i_map_35;
      end
      6'b100100 : begin
        _zz_shift_i_6_2 = shift_i_map_36;
      end
      6'b100101 : begin
        _zz_shift_i_6_2 = shift_i_map_37;
      end
      6'b100110 : begin
        _zz_shift_i_6_2 = shift_i_map_38;
      end
      default : begin
        _zz_shift_i_6_2 = shift_i_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_6_3)
      6'b000000 : begin
        _zz_shift_q_6_2 = shift_q_map_0;
      end
      6'b000001 : begin
        _zz_shift_q_6_2 = shift_q_map_1;
      end
      6'b000010 : begin
        _zz_shift_q_6_2 = shift_q_map_2;
      end
      6'b000011 : begin
        _zz_shift_q_6_2 = shift_q_map_3;
      end
      6'b000100 : begin
        _zz_shift_q_6_2 = shift_q_map_4;
      end
      6'b000101 : begin
        _zz_shift_q_6_2 = shift_q_map_5;
      end
      6'b000110 : begin
        _zz_shift_q_6_2 = shift_q_map_6;
      end
      6'b000111 : begin
        _zz_shift_q_6_2 = shift_q_map_7;
      end
      6'b001000 : begin
        _zz_shift_q_6_2 = shift_q_map_8;
      end
      6'b001001 : begin
        _zz_shift_q_6_2 = shift_q_map_9;
      end
      6'b001010 : begin
        _zz_shift_q_6_2 = shift_q_map_10;
      end
      6'b001011 : begin
        _zz_shift_q_6_2 = shift_q_map_11;
      end
      6'b001100 : begin
        _zz_shift_q_6_2 = shift_q_map_12;
      end
      6'b001101 : begin
        _zz_shift_q_6_2 = shift_q_map_13;
      end
      6'b001110 : begin
        _zz_shift_q_6_2 = shift_q_map_14;
      end
      6'b001111 : begin
        _zz_shift_q_6_2 = shift_q_map_15;
      end
      6'b010000 : begin
        _zz_shift_q_6_2 = shift_q_map_16;
      end
      6'b010001 : begin
        _zz_shift_q_6_2 = shift_q_map_17;
      end
      6'b010010 : begin
        _zz_shift_q_6_2 = shift_q_map_18;
      end
      6'b010011 : begin
        _zz_shift_q_6_2 = shift_q_map_19;
      end
      6'b010100 : begin
        _zz_shift_q_6_2 = shift_q_map_20;
      end
      6'b010101 : begin
        _zz_shift_q_6_2 = shift_q_map_21;
      end
      6'b010110 : begin
        _zz_shift_q_6_2 = shift_q_map_22;
      end
      6'b010111 : begin
        _zz_shift_q_6_2 = shift_q_map_23;
      end
      6'b011000 : begin
        _zz_shift_q_6_2 = shift_q_map_24;
      end
      6'b011001 : begin
        _zz_shift_q_6_2 = shift_q_map_25;
      end
      6'b011010 : begin
        _zz_shift_q_6_2 = shift_q_map_26;
      end
      6'b011011 : begin
        _zz_shift_q_6_2 = shift_q_map_27;
      end
      6'b011100 : begin
        _zz_shift_q_6_2 = shift_q_map_28;
      end
      6'b011101 : begin
        _zz_shift_q_6_2 = shift_q_map_29;
      end
      6'b011110 : begin
        _zz_shift_q_6_2 = shift_q_map_30;
      end
      6'b011111 : begin
        _zz_shift_q_6_2 = shift_q_map_31;
      end
      6'b100000 : begin
        _zz_shift_q_6_2 = shift_q_map_32;
      end
      6'b100001 : begin
        _zz_shift_q_6_2 = shift_q_map_33;
      end
      6'b100010 : begin
        _zz_shift_q_6_2 = shift_q_map_34;
      end
      6'b100011 : begin
        _zz_shift_q_6_2 = shift_q_map_35;
      end
      6'b100100 : begin
        _zz_shift_q_6_2 = shift_q_map_36;
      end
      6'b100101 : begin
        _zz_shift_q_6_2 = shift_q_map_37;
      end
      6'b100110 : begin
        _zz_shift_q_6_2 = shift_q_map_38;
      end
      default : begin
        _zz_shift_q_6_2 = shift_q_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_7_3)
      6'b000000 : begin
        _zz_shift_i_7_2 = shift_i_map_0;
      end
      6'b000001 : begin
        _zz_shift_i_7_2 = shift_i_map_1;
      end
      6'b000010 : begin
        _zz_shift_i_7_2 = shift_i_map_2;
      end
      6'b000011 : begin
        _zz_shift_i_7_2 = shift_i_map_3;
      end
      6'b000100 : begin
        _zz_shift_i_7_2 = shift_i_map_4;
      end
      6'b000101 : begin
        _zz_shift_i_7_2 = shift_i_map_5;
      end
      6'b000110 : begin
        _zz_shift_i_7_2 = shift_i_map_6;
      end
      6'b000111 : begin
        _zz_shift_i_7_2 = shift_i_map_7;
      end
      6'b001000 : begin
        _zz_shift_i_7_2 = shift_i_map_8;
      end
      6'b001001 : begin
        _zz_shift_i_7_2 = shift_i_map_9;
      end
      6'b001010 : begin
        _zz_shift_i_7_2 = shift_i_map_10;
      end
      6'b001011 : begin
        _zz_shift_i_7_2 = shift_i_map_11;
      end
      6'b001100 : begin
        _zz_shift_i_7_2 = shift_i_map_12;
      end
      6'b001101 : begin
        _zz_shift_i_7_2 = shift_i_map_13;
      end
      6'b001110 : begin
        _zz_shift_i_7_2 = shift_i_map_14;
      end
      6'b001111 : begin
        _zz_shift_i_7_2 = shift_i_map_15;
      end
      6'b010000 : begin
        _zz_shift_i_7_2 = shift_i_map_16;
      end
      6'b010001 : begin
        _zz_shift_i_7_2 = shift_i_map_17;
      end
      6'b010010 : begin
        _zz_shift_i_7_2 = shift_i_map_18;
      end
      6'b010011 : begin
        _zz_shift_i_7_2 = shift_i_map_19;
      end
      6'b010100 : begin
        _zz_shift_i_7_2 = shift_i_map_20;
      end
      6'b010101 : begin
        _zz_shift_i_7_2 = shift_i_map_21;
      end
      6'b010110 : begin
        _zz_shift_i_7_2 = shift_i_map_22;
      end
      6'b010111 : begin
        _zz_shift_i_7_2 = shift_i_map_23;
      end
      6'b011000 : begin
        _zz_shift_i_7_2 = shift_i_map_24;
      end
      6'b011001 : begin
        _zz_shift_i_7_2 = shift_i_map_25;
      end
      6'b011010 : begin
        _zz_shift_i_7_2 = shift_i_map_26;
      end
      6'b011011 : begin
        _zz_shift_i_7_2 = shift_i_map_27;
      end
      6'b011100 : begin
        _zz_shift_i_7_2 = shift_i_map_28;
      end
      6'b011101 : begin
        _zz_shift_i_7_2 = shift_i_map_29;
      end
      6'b011110 : begin
        _zz_shift_i_7_2 = shift_i_map_30;
      end
      6'b011111 : begin
        _zz_shift_i_7_2 = shift_i_map_31;
      end
      6'b100000 : begin
        _zz_shift_i_7_2 = shift_i_map_32;
      end
      6'b100001 : begin
        _zz_shift_i_7_2 = shift_i_map_33;
      end
      6'b100010 : begin
        _zz_shift_i_7_2 = shift_i_map_34;
      end
      6'b100011 : begin
        _zz_shift_i_7_2 = shift_i_map_35;
      end
      6'b100100 : begin
        _zz_shift_i_7_2 = shift_i_map_36;
      end
      6'b100101 : begin
        _zz_shift_i_7_2 = shift_i_map_37;
      end
      6'b100110 : begin
        _zz_shift_i_7_2 = shift_i_map_38;
      end
      default : begin
        _zz_shift_i_7_2 = shift_i_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_7_3)
      6'b000000 : begin
        _zz_shift_q_7_2 = shift_q_map_0;
      end
      6'b000001 : begin
        _zz_shift_q_7_2 = shift_q_map_1;
      end
      6'b000010 : begin
        _zz_shift_q_7_2 = shift_q_map_2;
      end
      6'b000011 : begin
        _zz_shift_q_7_2 = shift_q_map_3;
      end
      6'b000100 : begin
        _zz_shift_q_7_2 = shift_q_map_4;
      end
      6'b000101 : begin
        _zz_shift_q_7_2 = shift_q_map_5;
      end
      6'b000110 : begin
        _zz_shift_q_7_2 = shift_q_map_6;
      end
      6'b000111 : begin
        _zz_shift_q_7_2 = shift_q_map_7;
      end
      6'b001000 : begin
        _zz_shift_q_7_2 = shift_q_map_8;
      end
      6'b001001 : begin
        _zz_shift_q_7_2 = shift_q_map_9;
      end
      6'b001010 : begin
        _zz_shift_q_7_2 = shift_q_map_10;
      end
      6'b001011 : begin
        _zz_shift_q_7_2 = shift_q_map_11;
      end
      6'b001100 : begin
        _zz_shift_q_7_2 = shift_q_map_12;
      end
      6'b001101 : begin
        _zz_shift_q_7_2 = shift_q_map_13;
      end
      6'b001110 : begin
        _zz_shift_q_7_2 = shift_q_map_14;
      end
      6'b001111 : begin
        _zz_shift_q_7_2 = shift_q_map_15;
      end
      6'b010000 : begin
        _zz_shift_q_7_2 = shift_q_map_16;
      end
      6'b010001 : begin
        _zz_shift_q_7_2 = shift_q_map_17;
      end
      6'b010010 : begin
        _zz_shift_q_7_2 = shift_q_map_18;
      end
      6'b010011 : begin
        _zz_shift_q_7_2 = shift_q_map_19;
      end
      6'b010100 : begin
        _zz_shift_q_7_2 = shift_q_map_20;
      end
      6'b010101 : begin
        _zz_shift_q_7_2 = shift_q_map_21;
      end
      6'b010110 : begin
        _zz_shift_q_7_2 = shift_q_map_22;
      end
      6'b010111 : begin
        _zz_shift_q_7_2 = shift_q_map_23;
      end
      6'b011000 : begin
        _zz_shift_q_7_2 = shift_q_map_24;
      end
      6'b011001 : begin
        _zz_shift_q_7_2 = shift_q_map_25;
      end
      6'b011010 : begin
        _zz_shift_q_7_2 = shift_q_map_26;
      end
      6'b011011 : begin
        _zz_shift_q_7_2 = shift_q_map_27;
      end
      6'b011100 : begin
        _zz_shift_q_7_2 = shift_q_map_28;
      end
      6'b011101 : begin
        _zz_shift_q_7_2 = shift_q_map_29;
      end
      6'b011110 : begin
        _zz_shift_q_7_2 = shift_q_map_30;
      end
      6'b011111 : begin
        _zz_shift_q_7_2 = shift_q_map_31;
      end
      6'b100000 : begin
        _zz_shift_q_7_2 = shift_q_map_32;
      end
      6'b100001 : begin
        _zz_shift_q_7_2 = shift_q_map_33;
      end
      6'b100010 : begin
        _zz_shift_q_7_2 = shift_q_map_34;
      end
      6'b100011 : begin
        _zz_shift_q_7_2 = shift_q_map_35;
      end
      6'b100100 : begin
        _zz_shift_q_7_2 = shift_q_map_36;
      end
      6'b100101 : begin
        _zz_shift_q_7_2 = shift_q_map_37;
      end
      6'b100110 : begin
        _zz_shift_q_7_2 = shift_q_map_38;
      end
      default : begin
        _zz_shift_q_7_2 = shift_q_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_0_5)
      6'b000000 : begin
        _zz_shift_i_0_4 = shift_i_map_0;
      end
      6'b000001 : begin
        _zz_shift_i_0_4 = shift_i_map_1;
      end
      6'b000010 : begin
        _zz_shift_i_0_4 = shift_i_map_2;
      end
      6'b000011 : begin
        _zz_shift_i_0_4 = shift_i_map_3;
      end
      6'b000100 : begin
        _zz_shift_i_0_4 = shift_i_map_4;
      end
      6'b000101 : begin
        _zz_shift_i_0_4 = shift_i_map_5;
      end
      6'b000110 : begin
        _zz_shift_i_0_4 = shift_i_map_6;
      end
      6'b000111 : begin
        _zz_shift_i_0_4 = shift_i_map_7;
      end
      6'b001000 : begin
        _zz_shift_i_0_4 = shift_i_map_8;
      end
      6'b001001 : begin
        _zz_shift_i_0_4 = shift_i_map_9;
      end
      6'b001010 : begin
        _zz_shift_i_0_4 = shift_i_map_10;
      end
      6'b001011 : begin
        _zz_shift_i_0_4 = shift_i_map_11;
      end
      6'b001100 : begin
        _zz_shift_i_0_4 = shift_i_map_12;
      end
      6'b001101 : begin
        _zz_shift_i_0_4 = shift_i_map_13;
      end
      6'b001110 : begin
        _zz_shift_i_0_4 = shift_i_map_14;
      end
      6'b001111 : begin
        _zz_shift_i_0_4 = shift_i_map_15;
      end
      6'b010000 : begin
        _zz_shift_i_0_4 = shift_i_map_16;
      end
      6'b010001 : begin
        _zz_shift_i_0_4 = shift_i_map_17;
      end
      6'b010010 : begin
        _zz_shift_i_0_4 = shift_i_map_18;
      end
      6'b010011 : begin
        _zz_shift_i_0_4 = shift_i_map_19;
      end
      6'b010100 : begin
        _zz_shift_i_0_4 = shift_i_map_20;
      end
      6'b010101 : begin
        _zz_shift_i_0_4 = shift_i_map_21;
      end
      6'b010110 : begin
        _zz_shift_i_0_4 = shift_i_map_22;
      end
      6'b010111 : begin
        _zz_shift_i_0_4 = shift_i_map_23;
      end
      6'b011000 : begin
        _zz_shift_i_0_4 = shift_i_map_24;
      end
      6'b011001 : begin
        _zz_shift_i_0_4 = shift_i_map_25;
      end
      6'b011010 : begin
        _zz_shift_i_0_4 = shift_i_map_26;
      end
      6'b011011 : begin
        _zz_shift_i_0_4 = shift_i_map_27;
      end
      6'b011100 : begin
        _zz_shift_i_0_4 = shift_i_map_28;
      end
      6'b011101 : begin
        _zz_shift_i_0_4 = shift_i_map_29;
      end
      6'b011110 : begin
        _zz_shift_i_0_4 = shift_i_map_30;
      end
      6'b011111 : begin
        _zz_shift_i_0_4 = shift_i_map_31;
      end
      6'b100000 : begin
        _zz_shift_i_0_4 = shift_i_map_32;
      end
      6'b100001 : begin
        _zz_shift_i_0_4 = shift_i_map_33;
      end
      6'b100010 : begin
        _zz_shift_i_0_4 = shift_i_map_34;
      end
      6'b100011 : begin
        _zz_shift_i_0_4 = shift_i_map_35;
      end
      6'b100100 : begin
        _zz_shift_i_0_4 = shift_i_map_36;
      end
      6'b100101 : begin
        _zz_shift_i_0_4 = shift_i_map_37;
      end
      6'b100110 : begin
        _zz_shift_i_0_4 = shift_i_map_38;
      end
      default : begin
        _zz_shift_i_0_4 = shift_i_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_0_5)
      6'b000000 : begin
        _zz_shift_q_0_4 = shift_q_map_0;
      end
      6'b000001 : begin
        _zz_shift_q_0_4 = shift_q_map_1;
      end
      6'b000010 : begin
        _zz_shift_q_0_4 = shift_q_map_2;
      end
      6'b000011 : begin
        _zz_shift_q_0_4 = shift_q_map_3;
      end
      6'b000100 : begin
        _zz_shift_q_0_4 = shift_q_map_4;
      end
      6'b000101 : begin
        _zz_shift_q_0_4 = shift_q_map_5;
      end
      6'b000110 : begin
        _zz_shift_q_0_4 = shift_q_map_6;
      end
      6'b000111 : begin
        _zz_shift_q_0_4 = shift_q_map_7;
      end
      6'b001000 : begin
        _zz_shift_q_0_4 = shift_q_map_8;
      end
      6'b001001 : begin
        _zz_shift_q_0_4 = shift_q_map_9;
      end
      6'b001010 : begin
        _zz_shift_q_0_4 = shift_q_map_10;
      end
      6'b001011 : begin
        _zz_shift_q_0_4 = shift_q_map_11;
      end
      6'b001100 : begin
        _zz_shift_q_0_4 = shift_q_map_12;
      end
      6'b001101 : begin
        _zz_shift_q_0_4 = shift_q_map_13;
      end
      6'b001110 : begin
        _zz_shift_q_0_4 = shift_q_map_14;
      end
      6'b001111 : begin
        _zz_shift_q_0_4 = shift_q_map_15;
      end
      6'b010000 : begin
        _zz_shift_q_0_4 = shift_q_map_16;
      end
      6'b010001 : begin
        _zz_shift_q_0_4 = shift_q_map_17;
      end
      6'b010010 : begin
        _zz_shift_q_0_4 = shift_q_map_18;
      end
      6'b010011 : begin
        _zz_shift_q_0_4 = shift_q_map_19;
      end
      6'b010100 : begin
        _zz_shift_q_0_4 = shift_q_map_20;
      end
      6'b010101 : begin
        _zz_shift_q_0_4 = shift_q_map_21;
      end
      6'b010110 : begin
        _zz_shift_q_0_4 = shift_q_map_22;
      end
      6'b010111 : begin
        _zz_shift_q_0_4 = shift_q_map_23;
      end
      6'b011000 : begin
        _zz_shift_q_0_4 = shift_q_map_24;
      end
      6'b011001 : begin
        _zz_shift_q_0_4 = shift_q_map_25;
      end
      6'b011010 : begin
        _zz_shift_q_0_4 = shift_q_map_26;
      end
      6'b011011 : begin
        _zz_shift_q_0_4 = shift_q_map_27;
      end
      6'b011100 : begin
        _zz_shift_q_0_4 = shift_q_map_28;
      end
      6'b011101 : begin
        _zz_shift_q_0_4 = shift_q_map_29;
      end
      6'b011110 : begin
        _zz_shift_q_0_4 = shift_q_map_30;
      end
      6'b011111 : begin
        _zz_shift_q_0_4 = shift_q_map_31;
      end
      6'b100000 : begin
        _zz_shift_q_0_4 = shift_q_map_32;
      end
      6'b100001 : begin
        _zz_shift_q_0_4 = shift_q_map_33;
      end
      6'b100010 : begin
        _zz_shift_q_0_4 = shift_q_map_34;
      end
      6'b100011 : begin
        _zz_shift_q_0_4 = shift_q_map_35;
      end
      6'b100100 : begin
        _zz_shift_q_0_4 = shift_q_map_36;
      end
      6'b100101 : begin
        _zz_shift_q_0_4 = shift_q_map_37;
      end
      6'b100110 : begin
        _zz_shift_q_0_4 = shift_q_map_38;
      end
      default : begin
        _zz_shift_q_0_4 = shift_q_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_1_5)
      6'b000000 : begin
        _zz_shift_i_1_4 = shift_i_map_0;
      end
      6'b000001 : begin
        _zz_shift_i_1_4 = shift_i_map_1;
      end
      6'b000010 : begin
        _zz_shift_i_1_4 = shift_i_map_2;
      end
      6'b000011 : begin
        _zz_shift_i_1_4 = shift_i_map_3;
      end
      6'b000100 : begin
        _zz_shift_i_1_4 = shift_i_map_4;
      end
      6'b000101 : begin
        _zz_shift_i_1_4 = shift_i_map_5;
      end
      6'b000110 : begin
        _zz_shift_i_1_4 = shift_i_map_6;
      end
      6'b000111 : begin
        _zz_shift_i_1_4 = shift_i_map_7;
      end
      6'b001000 : begin
        _zz_shift_i_1_4 = shift_i_map_8;
      end
      6'b001001 : begin
        _zz_shift_i_1_4 = shift_i_map_9;
      end
      6'b001010 : begin
        _zz_shift_i_1_4 = shift_i_map_10;
      end
      6'b001011 : begin
        _zz_shift_i_1_4 = shift_i_map_11;
      end
      6'b001100 : begin
        _zz_shift_i_1_4 = shift_i_map_12;
      end
      6'b001101 : begin
        _zz_shift_i_1_4 = shift_i_map_13;
      end
      6'b001110 : begin
        _zz_shift_i_1_4 = shift_i_map_14;
      end
      6'b001111 : begin
        _zz_shift_i_1_4 = shift_i_map_15;
      end
      6'b010000 : begin
        _zz_shift_i_1_4 = shift_i_map_16;
      end
      6'b010001 : begin
        _zz_shift_i_1_4 = shift_i_map_17;
      end
      6'b010010 : begin
        _zz_shift_i_1_4 = shift_i_map_18;
      end
      6'b010011 : begin
        _zz_shift_i_1_4 = shift_i_map_19;
      end
      6'b010100 : begin
        _zz_shift_i_1_4 = shift_i_map_20;
      end
      6'b010101 : begin
        _zz_shift_i_1_4 = shift_i_map_21;
      end
      6'b010110 : begin
        _zz_shift_i_1_4 = shift_i_map_22;
      end
      6'b010111 : begin
        _zz_shift_i_1_4 = shift_i_map_23;
      end
      6'b011000 : begin
        _zz_shift_i_1_4 = shift_i_map_24;
      end
      6'b011001 : begin
        _zz_shift_i_1_4 = shift_i_map_25;
      end
      6'b011010 : begin
        _zz_shift_i_1_4 = shift_i_map_26;
      end
      6'b011011 : begin
        _zz_shift_i_1_4 = shift_i_map_27;
      end
      6'b011100 : begin
        _zz_shift_i_1_4 = shift_i_map_28;
      end
      6'b011101 : begin
        _zz_shift_i_1_4 = shift_i_map_29;
      end
      6'b011110 : begin
        _zz_shift_i_1_4 = shift_i_map_30;
      end
      6'b011111 : begin
        _zz_shift_i_1_4 = shift_i_map_31;
      end
      6'b100000 : begin
        _zz_shift_i_1_4 = shift_i_map_32;
      end
      6'b100001 : begin
        _zz_shift_i_1_4 = shift_i_map_33;
      end
      6'b100010 : begin
        _zz_shift_i_1_4 = shift_i_map_34;
      end
      6'b100011 : begin
        _zz_shift_i_1_4 = shift_i_map_35;
      end
      6'b100100 : begin
        _zz_shift_i_1_4 = shift_i_map_36;
      end
      6'b100101 : begin
        _zz_shift_i_1_4 = shift_i_map_37;
      end
      6'b100110 : begin
        _zz_shift_i_1_4 = shift_i_map_38;
      end
      default : begin
        _zz_shift_i_1_4 = shift_i_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_1_5)
      6'b000000 : begin
        _zz_shift_q_1_4 = shift_q_map_0;
      end
      6'b000001 : begin
        _zz_shift_q_1_4 = shift_q_map_1;
      end
      6'b000010 : begin
        _zz_shift_q_1_4 = shift_q_map_2;
      end
      6'b000011 : begin
        _zz_shift_q_1_4 = shift_q_map_3;
      end
      6'b000100 : begin
        _zz_shift_q_1_4 = shift_q_map_4;
      end
      6'b000101 : begin
        _zz_shift_q_1_4 = shift_q_map_5;
      end
      6'b000110 : begin
        _zz_shift_q_1_4 = shift_q_map_6;
      end
      6'b000111 : begin
        _zz_shift_q_1_4 = shift_q_map_7;
      end
      6'b001000 : begin
        _zz_shift_q_1_4 = shift_q_map_8;
      end
      6'b001001 : begin
        _zz_shift_q_1_4 = shift_q_map_9;
      end
      6'b001010 : begin
        _zz_shift_q_1_4 = shift_q_map_10;
      end
      6'b001011 : begin
        _zz_shift_q_1_4 = shift_q_map_11;
      end
      6'b001100 : begin
        _zz_shift_q_1_4 = shift_q_map_12;
      end
      6'b001101 : begin
        _zz_shift_q_1_4 = shift_q_map_13;
      end
      6'b001110 : begin
        _zz_shift_q_1_4 = shift_q_map_14;
      end
      6'b001111 : begin
        _zz_shift_q_1_4 = shift_q_map_15;
      end
      6'b010000 : begin
        _zz_shift_q_1_4 = shift_q_map_16;
      end
      6'b010001 : begin
        _zz_shift_q_1_4 = shift_q_map_17;
      end
      6'b010010 : begin
        _zz_shift_q_1_4 = shift_q_map_18;
      end
      6'b010011 : begin
        _zz_shift_q_1_4 = shift_q_map_19;
      end
      6'b010100 : begin
        _zz_shift_q_1_4 = shift_q_map_20;
      end
      6'b010101 : begin
        _zz_shift_q_1_4 = shift_q_map_21;
      end
      6'b010110 : begin
        _zz_shift_q_1_4 = shift_q_map_22;
      end
      6'b010111 : begin
        _zz_shift_q_1_4 = shift_q_map_23;
      end
      6'b011000 : begin
        _zz_shift_q_1_4 = shift_q_map_24;
      end
      6'b011001 : begin
        _zz_shift_q_1_4 = shift_q_map_25;
      end
      6'b011010 : begin
        _zz_shift_q_1_4 = shift_q_map_26;
      end
      6'b011011 : begin
        _zz_shift_q_1_4 = shift_q_map_27;
      end
      6'b011100 : begin
        _zz_shift_q_1_4 = shift_q_map_28;
      end
      6'b011101 : begin
        _zz_shift_q_1_4 = shift_q_map_29;
      end
      6'b011110 : begin
        _zz_shift_q_1_4 = shift_q_map_30;
      end
      6'b011111 : begin
        _zz_shift_q_1_4 = shift_q_map_31;
      end
      6'b100000 : begin
        _zz_shift_q_1_4 = shift_q_map_32;
      end
      6'b100001 : begin
        _zz_shift_q_1_4 = shift_q_map_33;
      end
      6'b100010 : begin
        _zz_shift_q_1_4 = shift_q_map_34;
      end
      6'b100011 : begin
        _zz_shift_q_1_4 = shift_q_map_35;
      end
      6'b100100 : begin
        _zz_shift_q_1_4 = shift_q_map_36;
      end
      6'b100101 : begin
        _zz_shift_q_1_4 = shift_q_map_37;
      end
      6'b100110 : begin
        _zz_shift_q_1_4 = shift_q_map_38;
      end
      default : begin
        _zz_shift_q_1_4 = shift_q_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_2_5)
      6'b000000 : begin
        _zz_shift_i_2_4 = shift_i_map_0;
      end
      6'b000001 : begin
        _zz_shift_i_2_4 = shift_i_map_1;
      end
      6'b000010 : begin
        _zz_shift_i_2_4 = shift_i_map_2;
      end
      6'b000011 : begin
        _zz_shift_i_2_4 = shift_i_map_3;
      end
      6'b000100 : begin
        _zz_shift_i_2_4 = shift_i_map_4;
      end
      6'b000101 : begin
        _zz_shift_i_2_4 = shift_i_map_5;
      end
      6'b000110 : begin
        _zz_shift_i_2_4 = shift_i_map_6;
      end
      6'b000111 : begin
        _zz_shift_i_2_4 = shift_i_map_7;
      end
      6'b001000 : begin
        _zz_shift_i_2_4 = shift_i_map_8;
      end
      6'b001001 : begin
        _zz_shift_i_2_4 = shift_i_map_9;
      end
      6'b001010 : begin
        _zz_shift_i_2_4 = shift_i_map_10;
      end
      6'b001011 : begin
        _zz_shift_i_2_4 = shift_i_map_11;
      end
      6'b001100 : begin
        _zz_shift_i_2_4 = shift_i_map_12;
      end
      6'b001101 : begin
        _zz_shift_i_2_4 = shift_i_map_13;
      end
      6'b001110 : begin
        _zz_shift_i_2_4 = shift_i_map_14;
      end
      6'b001111 : begin
        _zz_shift_i_2_4 = shift_i_map_15;
      end
      6'b010000 : begin
        _zz_shift_i_2_4 = shift_i_map_16;
      end
      6'b010001 : begin
        _zz_shift_i_2_4 = shift_i_map_17;
      end
      6'b010010 : begin
        _zz_shift_i_2_4 = shift_i_map_18;
      end
      6'b010011 : begin
        _zz_shift_i_2_4 = shift_i_map_19;
      end
      6'b010100 : begin
        _zz_shift_i_2_4 = shift_i_map_20;
      end
      6'b010101 : begin
        _zz_shift_i_2_4 = shift_i_map_21;
      end
      6'b010110 : begin
        _zz_shift_i_2_4 = shift_i_map_22;
      end
      6'b010111 : begin
        _zz_shift_i_2_4 = shift_i_map_23;
      end
      6'b011000 : begin
        _zz_shift_i_2_4 = shift_i_map_24;
      end
      6'b011001 : begin
        _zz_shift_i_2_4 = shift_i_map_25;
      end
      6'b011010 : begin
        _zz_shift_i_2_4 = shift_i_map_26;
      end
      6'b011011 : begin
        _zz_shift_i_2_4 = shift_i_map_27;
      end
      6'b011100 : begin
        _zz_shift_i_2_4 = shift_i_map_28;
      end
      6'b011101 : begin
        _zz_shift_i_2_4 = shift_i_map_29;
      end
      6'b011110 : begin
        _zz_shift_i_2_4 = shift_i_map_30;
      end
      6'b011111 : begin
        _zz_shift_i_2_4 = shift_i_map_31;
      end
      6'b100000 : begin
        _zz_shift_i_2_4 = shift_i_map_32;
      end
      6'b100001 : begin
        _zz_shift_i_2_4 = shift_i_map_33;
      end
      6'b100010 : begin
        _zz_shift_i_2_4 = shift_i_map_34;
      end
      6'b100011 : begin
        _zz_shift_i_2_4 = shift_i_map_35;
      end
      6'b100100 : begin
        _zz_shift_i_2_4 = shift_i_map_36;
      end
      6'b100101 : begin
        _zz_shift_i_2_4 = shift_i_map_37;
      end
      6'b100110 : begin
        _zz_shift_i_2_4 = shift_i_map_38;
      end
      default : begin
        _zz_shift_i_2_4 = shift_i_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_2_5)
      6'b000000 : begin
        _zz_shift_q_2_4 = shift_q_map_0;
      end
      6'b000001 : begin
        _zz_shift_q_2_4 = shift_q_map_1;
      end
      6'b000010 : begin
        _zz_shift_q_2_4 = shift_q_map_2;
      end
      6'b000011 : begin
        _zz_shift_q_2_4 = shift_q_map_3;
      end
      6'b000100 : begin
        _zz_shift_q_2_4 = shift_q_map_4;
      end
      6'b000101 : begin
        _zz_shift_q_2_4 = shift_q_map_5;
      end
      6'b000110 : begin
        _zz_shift_q_2_4 = shift_q_map_6;
      end
      6'b000111 : begin
        _zz_shift_q_2_4 = shift_q_map_7;
      end
      6'b001000 : begin
        _zz_shift_q_2_4 = shift_q_map_8;
      end
      6'b001001 : begin
        _zz_shift_q_2_4 = shift_q_map_9;
      end
      6'b001010 : begin
        _zz_shift_q_2_4 = shift_q_map_10;
      end
      6'b001011 : begin
        _zz_shift_q_2_4 = shift_q_map_11;
      end
      6'b001100 : begin
        _zz_shift_q_2_4 = shift_q_map_12;
      end
      6'b001101 : begin
        _zz_shift_q_2_4 = shift_q_map_13;
      end
      6'b001110 : begin
        _zz_shift_q_2_4 = shift_q_map_14;
      end
      6'b001111 : begin
        _zz_shift_q_2_4 = shift_q_map_15;
      end
      6'b010000 : begin
        _zz_shift_q_2_4 = shift_q_map_16;
      end
      6'b010001 : begin
        _zz_shift_q_2_4 = shift_q_map_17;
      end
      6'b010010 : begin
        _zz_shift_q_2_4 = shift_q_map_18;
      end
      6'b010011 : begin
        _zz_shift_q_2_4 = shift_q_map_19;
      end
      6'b010100 : begin
        _zz_shift_q_2_4 = shift_q_map_20;
      end
      6'b010101 : begin
        _zz_shift_q_2_4 = shift_q_map_21;
      end
      6'b010110 : begin
        _zz_shift_q_2_4 = shift_q_map_22;
      end
      6'b010111 : begin
        _zz_shift_q_2_4 = shift_q_map_23;
      end
      6'b011000 : begin
        _zz_shift_q_2_4 = shift_q_map_24;
      end
      6'b011001 : begin
        _zz_shift_q_2_4 = shift_q_map_25;
      end
      6'b011010 : begin
        _zz_shift_q_2_4 = shift_q_map_26;
      end
      6'b011011 : begin
        _zz_shift_q_2_4 = shift_q_map_27;
      end
      6'b011100 : begin
        _zz_shift_q_2_4 = shift_q_map_28;
      end
      6'b011101 : begin
        _zz_shift_q_2_4 = shift_q_map_29;
      end
      6'b011110 : begin
        _zz_shift_q_2_4 = shift_q_map_30;
      end
      6'b011111 : begin
        _zz_shift_q_2_4 = shift_q_map_31;
      end
      6'b100000 : begin
        _zz_shift_q_2_4 = shift_q_map_32;
      end
      6'b100001 : begin
        _zz_shift_q_2_4 = shift_q_map_33;
      end
      6'b100010 : begin
        _zz_shift_q_2_4 = shift_q_map_34;
      end
      6'b100011 : begin
        _zz_shift_q_2_4 = shift_q_map_35;
      end
      6'b100100 : begin
        _zz_shift_q_2_4 = shift_q_map_36;
      end
      6'b100101 : begin
        _zz_shift_q_2_4 = shift_q_map_37;
      end
      6'b100110 : begin
        _zz_shift_q_2_4 = shift_q_map_38;
      end
      default : begin
        _zz_shift_q_2_4 = shift_q_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_3_5)
      6'b000000 : begin
        _zz_shift_i_3_4 = shift_i_map_0;
      end
      6'b000001 : begin
        _zz_shift_i_3_4 = shift_i_map_1;
      end
      6'b000010 : begin
        _zz_shift_i_3_4 = shift_i_map_2;
      end
      6'b000011 : begin
        _zz_shift_i_3_4 = shift_i_map_3;
      end
      6'b000100 : begin
        _zz_shift_i_3_4 = shift_i_map_4;
      end
      6'b000101 : begin
        _zz_shift_i_3_4 = shift_i_map_5;
      end
      6'b000110 : begin
        _zz_shift_i_3_4 = shift_i_map_6;
      end
      6'b000111 : begin
        _zz_shift_i_3_4 = shift_i_map_7;
      end
      6'b001000 : begin
        _zz_shift_i_3_4 = shift_i_map_8;
      end
      6'b001001 : begin
        _zz_shift_i_3_4 = shift_i_map_9;
      end
      6'b001010 : begin
        _zz_shift_i_3_4 = shift_i_map_10;
      end
      6'b001011 : begin
        _zz_shift_i_3_4 = shift_i_map_11;
      end
      6'b001100 : begin
        _zz_shift_i_3_4 = shift_i_map_12;
      end
      6'b001101 : begin
        _zz_shift_i_3_4 = shift_i_map_13;
      end
      6'b001110 : begin
        _zz_shift_i_3_4 = shift_i_map_14;
      end
      6'b001111 : begin
        _zz_shift_i_3_4 = shift_i_map_15;
      end
      6'b010000 : begin
        _zz_shift_i_3_4 = shift_i_map_16;
      end
      6'b010001 : begin
        _zz_shift_i_3_4 = shift_i_map_17;
      end
      6'b010010 : begin
        _zz_shift_i_3_4 = shift_i_map_18;
      end
      6'b010011 : begin
        _zz_shift_i_3_4 = shift_i_map_19;
      end
      6'b010100 : begin
        _zz_shift_i_3_4 = shift_i_map_20;
      end
      6'b010101 : begin
        _zz_shift_i_3_4 = shift_i_map_21;
      end
      6'b010110 : begin
        _zz_shift_i_3_4 = shift_i_map_22;
      end
      6'b010111 : begin
        _zz_shift_i_3_4 = shift_i_map_23;
      end
      6'b011000 : begin
        _zz_shift_i_3_4 = shift_i_map_24;
      end
      6'b011001 : begin
        _zz_shift_i_3_4 = shift_i_map_25;
      end
      6'b011010 : begin
        _zz_shift_i_3_4 = shift_i_map_26;
      end
      6'b011011 : begin
        _zz_shift_i_3_4 = shift_i_map_27;
      end
      6'b011100 : begin
        _zz_shift_i_3_4 = shift_i_map_28;
      end
      6'b011101 : begin
        _zz_shift_i_3_4 = shift_i_map_29;
      end
      6'b011110 : begin
        _zz_shift_i_3_4 = shift_i_map_30;
      end
      6'b011111 : begin
        _zz_shift_i_3_4 = shift_i_map_31;
      end
      6'b100000 : begin
        _zz_shift_i_3_4 = shift_i_map_32;
      end
      6'b100001 : begin
        _zz_shift_i_3_4 = shift_i_map_33;
      end
      6'b100010 : begin
        _zz_shift_i_3_4 = shift_i_map_34;
      end
      6'b100011 : begin
        _zz_shift_i_3_4 = shift_i_map_35;
      end
      6'b100100 : begin
        _zz_shift_i_3_4 = shift_i_map_36;
      end
      6'b100101 : begin
        _zz_shift_i_3_4 = shift_i_map_37;
      end
      6'b100110 : begin
        _zz_shift_i_3_4 = shift_i_map_38;
      end
      default : begin
        _zz_shift_i_3_4 = shift_i_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_3_5)
      6'b000000 : begin
        _zz_shift_q_3_4 = shift_q_map_0;
      end
      6'b000001 : begin
        _zz_shift_q_3_4 = shift_q_map_1;
      end
      6'b000010 : begin
        _zz_shift_q_3_4 = shift_q_map_2;
      end
      6'b000011 : begin
        _zz_shift_q_3_4 = shift_q_map_3;
      end
      6'b000100 : begin
        _zz_shift_q_3_4 = shift_q_map_4;
      end
      6'b000101 : begin
        _zz_shift_q_3_4 = shift_q_map_5;
      end
      6'b000110 : begin
        _zz_shift_q_3_4 = shift_q_map_6;
      end
      6'b000111 : begin
        _zz_shift_q_3_4 = shift_q_map_7;
      end
      6'b001000 : begin
        _zz_shift_q_3_4 = shift_q_map_8;
      end
      6'b001001 : begin
        _zz_shift_q_3_4 = shift_q_map_9;
      end
      6'b001010 : begin
        _zz_shift_q_3_4 = shift_q_map_10;
      end
      6'b001011 : begin
        _zz_shift_q_3_4 = shift_q_map_11;
      end
      6'b001100 : begin
        _zz_shift_q_3_4 = shift_q_map_12;
      end
      6'b001101 : begin
        _zz_shift_q_3_4 = shift_q_map_13;
      end
      6'b001110 : begin
        _zz_shift_q_3_4 = shift_q_map_14;
      end
      6'b001111 : begin
        _zz_shift_q_3_4 = shift_q_map_15;
      end
      6'b010000 : begin
        _zz_shift_q_3_4 = shift_q_map_16;
      end
      6'b010001 : begin
        _zz_shift_q_3_4 = shift_q_map_17;
      end
      6'b010010 : begin
        _zz_shift_q_3_4 = shift_q_map_18;
      end
      6'b010011 : begin
        _zz_shift_q_3_4 = shift_q_map_19;
      end
      6'b010100 : begin
        _zz_shift_q_3_4 = shift_q_map_20;
      end
      6'b010101 : begin
        _zz_shift_q_3_4 = shift_q_map_21;
      end
      6'b010110 : begin
        _zz_shift_q_3_4 = shift_q_map_22;
      end
      6'b010111 : begin
        _zz_shift_q_3_4 = shift_q_map_23;
      end
      6'b011000 : begin
        _zz_shift_q_3_4 = shift_q_map_24;
      end
      6'b011001 : begin
        _zz_shift_q_3_4 = shift_q_map_25;
      end
      6'b011010 : begin
        _zz_shift_q_3_4 = shift_q_map_26;
      end
      6'b011011 : begin
        _zz_shift_q_3_4 = shift_q_map_27;
      end
      6'b011100 : begin
        _zz_shift_q_3_4 = shift_q_map_28;
      end
      6'b011101 : begin
        _zz_shift_q_3_4 = shift_q_map_29;
      end
      6'b011110 : begin
        _zz_shift_q_3_4 = shift_q_map_30;
      end
      6'b011111 : begin
        _zz_shift_q_3_4 = shift_q_map_31;
      end
      6'b100000 : begin
        _zz_shift_q_3_4 = shift_q_map_32;
      end
      6'b100001 : begin
        _zz_shift_q_3_4 = shift_q_map_33;
      end
      6'b100010 : begin
        _zz_shift_q_3_4 = shift_q_map_34;
      end
      6'b100011 : begin
        _zz_shift_q_3_4 = shift_q_map_35;
      end
      6'b100100 : begin
        _zz_shift_q_3_4 = shift_q_map_36;
      end
      6'b100101 : begin
        _zz_shift_q_3_4 = shift_q_map_37;
      end
      6'b100110 : begin
        _zz_shift_q_3_4 = shift_q_map_38;
      end
      default : begin
        _zz_shift_q_3_4 = shift_q_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_4_5)
      6'b000000 : begin
        _zz_shift_i_4_4 = shift_i_map_0;
      end
      6'b000001 : begin
        _zz_shift_i_4_4 = shift_i_map_1;
      end
      6'b000010 : begin
        _zz_shift_i_4_4 = shift_i_map_2;
      end
      6'b000011 : begin
        _zz_shift_i_4_4 = shift_i_map_3;
      end
      6'b000100 : begin
        _zz_shift_i_4_4 = shift_i_map_4;
      end
      6'b000101 : begin
        _zz_shift_i_4_4 = shift_i_map_5;
      end
      6'b000110 : begin
        _zz_shift_i_4_4 = shift_i_map_6;
      end
      6'b000111 : begin
        _zz_shift_i_4_4 = shift_i_map_7;
      end
      6'b001000 : begin
        _zz_shift_i_4_4 = shift_i_map_8;
      end
      6'b001001 : begin
        _zz_shift_i_4_4 = shift_i_map_9;
      end
      6'b001010 : begin
        _zz_shift_i_4_4 = shift_i_map_10;
      end
      6'b001011 : begin
        _zz_shift_i_4_4 = shift_i_map_11;
      end
      6'b001100 : begin
        _zz_shift_i_4_4 = shift_i_map_12;
      end
      6'b001101 : begin
        _zz_shift_i_4_4 = shift_i_map_13;
      end
      6'b001110 : begin
        _zz_shift_i_4_4 = shift_i_map_14;
      end
      6'b001111 : begin
        _zz_shift_i_4_4 = shift_i_map_15;
      end
      6'b010000 : begin
        _zz_shift_i_4_4 = shift_i_map_16;
      end
      6'b010001 : begin
        _zz_shift_i_4_4 = shift_i_map_17;
      end
      6'b010010 : begin
        _zz_shift_i_4_4 = shift_i_map_18;
      end
      6'b010011 : begin
        _zz_shift_i_4_4 = shift_i_map_19;
      end
      6'b010100 : begin
        _zz_shift_i_4_4 = shift_i_map_20;
      end
      6'b010101 : begin
        _zz_shift_i_4_4 = shift_i_map_21;
      end
      6'b010110 : begin
        _zz_shift_i_4_4 = shift_i_map_22;
      end
      6'b010111 : begin
        _zz_shift_i_4_4 = shift_i_map_23;
      end
      6'b011000 : begin
        _zz_shift_i_4_4 = shift_i_map_24;
      end
      6'b011001 : begin
        _zz_shift_i_4_4 = shift_i_map_25;
      end
      6'b011010 : begin
        _zz_shift_i_4_4 = shift_i_map_26;
      end
      6'b011011 : begin
        _zz_shift_i_4_4 = shift_i_map_27;
      end
      6'b011100 : begin
        _zz_shift_i_4_4 = shift_i_map_28;
      end
      6'b011101 : begin
        _zz_shift_i_4_4 = shift_i_map_29;
      end
      6'b011110 : begin
        _zz_shift_i_4_4 = shift_i_map_30;
      end
      6'b011111 : begin
        _zz_shift_i_4_4 = shift_i_map_31;
      end
      6'b100000 : begin
        _zz_shift_i_4_4 = shift_i_map_32;
      end
      6'b100001 : begin
        _zz_shift_i_4_4 = shift_i_map_33;
      end
      6'b100010 : begin
        _zz_shift_i_4_4 = shift_i_map_34;
      end
      6'b100011 : begin
        _zz_shift_i_4_4 = shift_i_map_35;
      end
      6'b100100 : begin
        _zz_shift_i_4_4 = shift_i_map_36;
      end
      6'b100101 : begin
        _zz_shift_i_4_4 = shift_i_map_37;
      end
      6'b100110 : begin
        _zz_shift_i_4_4 = shift_i_map_38;
      end
      default : begin
        _zz_shift_i_4_4 = shift_i_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_4_5)
      6'b000000 : begin
        _zz_shift_q_4_4 = shift_q_map_0;
      end
      6'b000001 : begin
        _zz_shift_q_4_4 = shift_q_map_1;
      end
      6'b000010 : begin
        _zz_shift_q_4_4 = shift_q_map_2;
      end
      6'b000011 : begin
        _zz_shift_q_4_4 = shift_q_map_3;
      end
      6'b000100 : begin
        _zz_shift_q_4_4 = shift_q_map_4;
      end
      6'b000101 : begin
        _zz_shift_q_4_4 = shift_q_map_5;
      end
      6'b000110 : begin
        _zz_shift_q_4_4 = shift_q_map_6;
      end
      6'b000111 : begin
        _zz_shift_q_4_4 = shift_q_map_7;
      end
      6'b001000 : begin
        _zz_shift_q_4_4 = shift_q_map_8;
      end
      6'b001001 : begin
        _zz_shift_q_4_4 = shift_q_map_9;
      end
      6'b001010 : begin
        _zz_shift_q_4_4 = shift_q_map_10;
      end
      6'b001011 : begin
        _zz_shift_q_4_4 = shift_q_map_11;
      end
      6'b001100 : begin
        _zz_shift_q_4_4 = shift_q_map_12;
      end
      6'b001101 : begin
        _zz_shift_q_4_4 = shift_q_map_13;
      end
      6'b001110 : begin
        _zz_shift_q_4_4 = shift_q_map_14;
      end
      6'b001111 : begin
        _zz_shift_q_4_4 = shift_q_map_15;
      end
      6'b010000 : begin
        _zz_shift_q_4_4 = shift_q_map_16;
      end
      6'b010001 : begin
        _zz_shift_q_4_4 = shift_q_map_17;
      end
      6'b010010 : begin
        _zz_shift_q_4_4 = shift_q_map_18;
      end
      6'b010011 : begin
        _zz_shift_q_4_4 = shift_q_map_19;
      end
      6'b010100 : begin
        _zz_shift_q_4_4 = shift_q_map_20;
      end
      6'b010101 : begin
        _zz_shift_q_4_4 = shift_q_map_21;
      end
      6'b010110 : begin
        _zz_shift_q_4_4 = shift_q_map_22;
      end
      6'b010111 : begin
        _zz_shift_q_4_4 = shift_q_map_23;
      end
      6'b011000 : begin
        _zz_shift_q_4_4 = shift_q_map_24;
      end
      6'b011001 : begin
        _zz_shift_q_4_4 = shift_q_map_25;
      end
      6'b011010 : begin
        _zz_shift_q_4_4 = shift_q_map_26;
      end
      6'b011011 : begin
        _zz_shift_q_4_4 = shift_q_map_27;
      end
      6'b011100 : begin
        _zz_shift_q_4_4 = shift_q_map_28;
      end
      6'b011101 : begin
        _zz_shift_q_4_4 = shift_q_map_29;
      end
      6'b011110 : begin
        _zz_shift_q_4_4 = shift_q_map_30;
      end
      6'b011111 : begin
        _zz_shift_q_4_4 = shift_q_map_31;
      end
      6'b100000 : begin
        _zz_shift_q_4_4 = shift_q_map_32;
      end
      6'b100001 : begin
        _zz_shift_q_4_4 = shift_q_map_33;
      end
      6'b100010 : begin
        _zz_shift_q_4_4 = shift_q_map_34;
      end
      6'b100011 : begin
        _zz_shift_q_4_4 = shift_q_map_35;
      end
      6'b100100 : begin
        _zz_shift_q_4_4 = shift_q_map_36;
      end
      6'b100101 : begin
        _zz_shift_q_4_4 = shift_q_map_37;
      end
      6'b100110 : begin
        _zz_shift_q_4_4 = shift_q_map_38;
      end
      default : begin
        _zz_shift_q_4_4 = shift_q_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_5_5)
      6'b000000 : begin
        _zz_shift_i_5_4 = shift_i_map_0;
      end
      6'b000001 : begin
        _zz_shift_i_5_4 = shift_i_map_1;
      end
      6'b000010 : begin
        _zz_shift_i_5_4 = shift_i_map_2;
      end
      6'b000011 : begin
        _zz_shift_i_5_4 = shift_i_map_3;
      end
      6'b000100 : begin
        _zz_shift_i_5_4 = shift_i_map_4;
      end
      6'b000101 : begin
        _zz_shift_i_5_4 = shift_i_map_5;
      end
      6'b000110 : begin
        _zz_shift_i_5_4 = shift_i_map_6;
      end
      6'b000111 : begin
        _zz_shift_i_5_4 = shift_i_map_7;
      end
      6'b001000 : begin
        _zz_shift_i_5_4 = shift_i_map_8;
      end
      6'b001001 : begin
        _zz_shift_i_5_4 = shift_i_map_9;
      end
      6'b001010 : begin
        _zz_shift_i_5_4 = shift_i_map_10;
      end
      6'b001011 : begin
        _zz_shift_i_5_4 = shift_i_map_11;
      end
      6'b001100 : begin
        _zz_shift_i_5_4 = shift_i_map_12;
      end
      6'b001101 : begin
        _zz_shift_i_5_4 = shift_i_map_13;
      end
      6'b001110 : begin
        _zz_shift_i_5_4 = shift_i_map_14;
      end
      6'b001111 : begin
        _zz_shift_i_5_4 = shift_i_map_15;
      end
      6'b010000 : begin
        _zz_shift_i_5_4 = shift_i_map_16;
      end
      6'b010001 : begin
        _zz_shift_i_5_4 = shift_i_map_17;
      end
      6'b010010 : begin
        _zz_shift_i_5_4 = shift_i_map_18;
      end
      6'b010011 : begin
        _zz_shift_i_5_4 = shift_i_map_19;
      end
      6'b010100 : begin
        _zz_shift_i_5_4 = shift_i_map_20;
      end
      6'b010101 : begin
        _zz_shift_i_5_4 = shift_i_map_21;
      end
      6'b010110 : begin
        _zz_shift_i_5_4 = shift_i_map_22;
      end
      6'b010111 : begin
        _zz_shift_i_5_4 = shift_i_map_23;
      end
      6'b011000 : begin
        _zz_shift_i_5_4 = shift_i_map_24;
      end
      6'b011001 : begin
        _zz_shift_i_5_4 = shift_i_map_25;
      end
      6'b011010 : begin
        _zz_shift_i_5_4 = shift_i_map_26;
      end
      6'b011011 : begin
        _zz_shift_i_5_4 = shift_i_map_27;
      end
      6'b011100 : begin
        _zz_shift_i_5_4 = shift_i_map_28;
      end
      6'b011101 : begin
        _zz_shift_i_5_4 = shift_i_map_29;
      end
      6'b011110 : begin
        _zz_shift_i_5_4 = shift_i_map_30;
      end
      6'b011111 : begin
        _zz_shift_i_5_4 = shift_i_map_31;
      end
      6'b100000 : begin
        _zz_shift_i_5_4 = shift_i_map_32;
      end
      6'b100001 : begin
        _zz_shift_i_5_4 = shift_i_map_33;
      end
      6'b100010 : begin
        _zz_shift_i_5_4 = shift_i_map_34;
      end
      6'b100011 : begin
        _zz_shift_i_5_4 = shift_i_map_35;
      end
      6'b100100 : begin
        _zz_shift_i_5_4 = shift_i_map_36;
      end
      6'b100101 : begin
        _zz_shift_i_5_4 = shift_i_map_37;
      end
      6'b100110 : begin
        _zz_shift_i_5_4 = shift_i_map_38;
      end
      default : begin
        _zz_shift_i_5_4 = shift_i_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_5_5)
      6'b000000 : begin
        _zz_shift_q_5_4 = shift_q_map_0;
      end
      6'b000001 : begin
        _zz_shift_q_5_4 = shift_q_map_1;
      end
      6'b000010 : begin
        _zz_shift_q_5_4 = shift_q_map_2;
      end
      6'b000011 : begin
        _zz_shift_q_5_4 = shift_q_map_3;
      end
      6'b000100 : begin
        _zz_shift_q_5_4 = shift_q_map_4;
      end
      6'b000101 : begin
        _zz_shift_q_5_4 = shift_q_map_5;
      end
      6'b000110 : begin
        _zz_shift_q_5_4 = shift_q_map_6;
      end
      6'b000111 : begin
        _zz_shift_q_5_4 = shift_q_map_7;
      end
      6'b001000 : begin
        _zz_shift_q_5_4 = shift_q_map_8;
      end
      6'b001001 : begin
        _zz_shift_q_5_4 = shift_q_map_9;
      end
      6'b001010 : begin
        _zz_shift_q_5_4 = shift_q_map_10;
      end
      6'b001011 : begin
        _zz_shift_q_5_4 = shift_q_map_11;
      end
      6'b001100 : begin
        _zz_shift_q_5_4 = shift_q_map_12;
      end
      6'b001101 : begin
        _zz_shift_q_5_4 = shift_q_map_13;
      end
      6'b001110 : begin
        _zz_shift_q_5_4 = shift_q_map_14;
      end
      6'b001111 : begin
        _zz_shift_q_5_4 = shift_q_map_15;
      end
      6'b010000 : begin
        _zz_shift_q_5_4 = shift_q_map_16;
      end
      6'b010001 : begin
        _zz_shift_q_5_4 = shift_q_map_17;
      end
      6'b010010 : begin
        _zz_shift_q_5_4 = shift_q_map_18;
      end
      6'b010011 : begin
        _zz_shift_q_5_4 = shift_q_map_19;
      end
      6'b010100 : begin
        _zz_shift_q_5_4 = shift_q_map_20;
      end
      6'b010101 : begin
        _zz_shift_q_5_4 = shift_q_map_21;
      end
      6'b010110 : begin
        _zz_shift_q_5_4 = shift_q_map_22;
      end
      6'b010111 : begin
        _zz_shift_q_5_4 = shift_q_map_23;
      end
      6'b011000 : begin
        _zz_shift_q_5_4 = shift_q_map_24;
      end
      6'b011001 : begin
        _zz_shift_q_5_4 = shift_q_map_25;
      end
      6'b011010 : begin
        _zz_shift_q_5_4 = shift_q_map_26;
      end
      6'b011011 : begin
        _zz_shift_q_5_4 = shift_q_map_27;
      end
      6'b011100 : begin
        _zz_shift_q_5_4 = shift_q_map_28;
      end
      6'b011101 : begin
        _zz_shift_q_5_4 = shift_q_map_29;
      end
      6'b011110 : begin
        _zz_shift_q_5_4 = shift_q_map_30;
      end
      6'b011111 : begin
        _zz_shift_q_5_4 = shift_q_map_31;
      end
      6'b100000 : begin
        _zz_shift_q_5_4 = shift_q_map_32;
      end
      6'b100001 : begin
        _zz_shift_q_5_4 = shift_q_map_33;
      end
      6'b100010 : begin
        _zz_shift_q_5_4 = shift_q_map_34;
      end
      6'b100011 : begin
        _zz_shift_q_5_4 = shift_q_map_35;
      end
      6'b100100 : begin
        _zz_shift_q_5_4 = shift_q_map_36;
      end
      6'b100101 : begin
        _zz_shift_q_5_4 = shift_q_map_37;
      end
      6'b100110 : begin
        _zz_shift_q_5_4 = shift_q_map_38;
      end
      default : begin
        _zz_shift_q_5_4 = shift_q_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_6_5)
      6'b000000 : begin
        _zz_shift_i_6_4 = shift_i_map_0;
      end
      6'b000001 : begin
        _zz_shift_i_6_4 = shift_i_map_1;
      end
      6'b000010 : begin
        _zz_shift_i_6_4 = shift_i_map_2;
      end
      6'b000011 : begin
        _zz_shift_i_6_4 = shift_i_map_3;
      end
      6'b000100 : begin
        _zz_shift_i_6_4 = shift_i_map_4;
      end
      6'b000101 : begin
        _zz_shift_i_6_4 = shift_i_map_5;
      end
      6'b000110 : begin
        _zz_shift_i_6_4 = shift_i_map_6;
      end
      6'b000111 : begin
        _zz_shift_i_6_4 = shift_i_map_7;
      end
      6'b001000 : begin
        _zz_shift_i_6_4 = shift_i_map_8;
      end
      6'b001001 : begin
        _zz_shift_i_6_4 = shift_i_map_9;
      end
      6'b001010 : begin
        _zz_shift_i_6_4 = shift_i_map_10;
      end
      6'b001011 : begin
        _zz_shift_i_6_4 = shift_i_map_11;
      end
      6'b001100 : begin
        _zz_shift_i_6_4 = shift_i_map_12;
      end
      6'b001101 : begin
        _zz_shift_i_6_4 = shift_i_map_13;
      end
      6'b001110 : begin
        _zz_shift_i_6_4 = shift_i_map_14;
      end
      6'b001111 : begin
        _zz_shift_i_6_4 = shift_i_map_15;
      end
      6'b010000 : begin
        _zz_shift_i_6_4 = shift_i_map_16;
      end
      6'b010001 : begin
        _zz_shift_i_6_4 = shift_i_map_17;
      end
      6'b010010 : begin
        _zz_shift_i_6_4 = shift_i_map_18;
      end
      6'b010011 : begin
        _zz_shift_i_6_4 = shift_i_map_19;
      end
      6'b010100 : begin
        _zz_shift_i_6_4 = shift_i_map_20;
      end
      6'b010101 : begin
        _zz_shift_i_6_4 = shift_i_map_21;
      end
      6'b010110 : begin
        _zz_shift_i_6_4 = shift_i_map_22;
      end
      6'b010111 : begin
        _zz_shift_i_6_4 = shift_i_map_23;
      end
      6'b011000 : begin
        _zz_shift_i_6_4 = shift_i_map_24;
      end
      6'b011001 : begin
        _zz_shift_i_6_4 = shift_i_map_25;
      end
      6'b011010 : begin
        _zz_shift_i_6_4 = shift_i_map_26;
      end
      6'b011011 : begin
        _zz_shift_i_6_4 = shift_i_map_27;
      end
      6'b011100 : begin
        _zz_shift_i_6_4 = shift_i_map_28;
      end
      6'b011101 : begin
        _zz_shift_i_6_4 = shift_i_map_29;
      end
      6'b011110 : begin
        _zz_shift_i_6_4 = shift_i_map_30;
      end
      6'b011111 : begin
        _zz_shift_i_6_4 = shift_i_map_31;
      end
      6'b100000 : begin
        _zz_shift_i_6_4 = shift_i_map_32;
      end
      6'b100001 : begin
        _zz_shift_i_6_4 = shift_i_map_33;
      end
      6'b100010 : begin
        _zz_shift_i_6_4 = shift_i_map_34;
      end
      6'b100011 : begin
        _zz_shift_i_6_4 = shift_i_map_35;
      end
      6'b100100 : begin
        _zz_shift_i_6_4 = shift_i_map_36;
      end
      6'b100101 : begin
        _zz_shift_i_6_4 = shift_i_map_37;
      end
      6'b100110 : begin
        _zz_shift_i_6_4 = shift_i_map_38;
      end
      default : begin
        _zz_shift_i_6_4 = shift_i_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_6_5)
      6'b000000 : begin
        _zz_shift_q_6_4 = shift_q_map_0;
      end
      6'b000001 : begin
        _zz_shift_q_6_4 = shift_q_map_1;
      end
      6'b000010 : begin
        _zz_shift_q_6_4 = shift_q_map_2;
      end
      6'b000011 : begin
        _zz_shift_q_6_4 = shift_q_map_3;
      end
      6'b000100 : begin
        _zz_shift_q_6_4 = shift_q_map_4;
      end
      6'b000101 : begin
        _zz_shift_q_6_4 = shift_q_map_5;
      end
      6'b000110 : begin
        _zz_shift_q_6_4 = shift_q_map_6;
      end
      6'b000111 : begin
        _zz_shift_q_6_4 = shift_q_map_7;
      end
      6'b001000 : begin
        _zz_shift_q_6_4 = shift_q_map_8;
      end
      6'b001001 : begin
        _zz_shift_q_6_4 = shift_q_map_9;
      end
      6'b001010 : begin
        _zz_shift_q_6_4 = shift_q_map_10;
      end
      6'b001011 : begin
        _zz_shift_q_6_4 = shift_q_map_11;
      end
      6'b001100 : begin
        _zz_shift_q_6_4 = shift_q_map_12;
      end
      6'b001101 : begin
        _zz_shift_q_6_4 = shift_q_map_13;
      end
      6'b001110 : begin
        _zz_shift_q_6_4 = shift_q_map_14;
      end
      6'b001111 : begin
        _zz_shift_q_6_4 = shift_q_map_15;
      end
      6'b010000 : begin
        _zz_shift_q_6_4 = shift_q_map_16;
      end
      6'b010001 : begin
        _zz_shift_q_6_4 = shift_q_map_17;
      end
      6'b010010 : begin
        _zz_shift_q_6_4 = shift_q_map_18;
      end
      6'b010011 : begin
        _zz_shift_q_6_4 = shift_q_map_19;
      end
      6'b010100 : begin
        _zz_shift_q_6_4 = shift_q_map_20;
      end
      6'b010101 : begin
        _zz_shift_q_6_4 = shift_q_map_21;
      end
      6'b010110 : begin
        _zz_shift_q_6_4 = shift_q_map_22;
      end
      6'b010111 : begin
        _zz_shift_q_6_4 = shift_q_map_23;
      end
      6'b011000 : begin
        _zz_shift_q_6_4 = shift_q_map_24;
      end
      6'b011001 : begin
        _zz_shift_q_6_4 = shift_q_map_25;
      end
      6'b011010 : begin
        _zz_shift_q_6_4 = shift_q_map_26;
      end
      6'b011011 : begin
        _zz_shift_q_6_4 = shift_q_map_27;
      end
      6'b011100 : begin
        _zz_shift_q_6_4 = shift_q_map_28;
      end
      6'b011101 : begin
        _zz_shift_q_6_4 = shift_q_map_29;
      end
      6'b011110 : begin
        _zz_shift_q_6_4 = shift_q_map_30;
      end
      6'b011111 : begin
        _zz_shift_q_6_4 = shift_q_map_31;
      end
      6'b100000 : begin
        _zz_shift_q_6_4 = shift_q_map_32;
      end
      6'b100001 : begin
        _zz_shift_q_6_4 = shift_q_map_33;
      end
      6'b100010 : begin
        _zz_shift_q_6_4 = shift_q_map_34;
      end
      6'b100011 : begin
        _zz_shift_q_6_4 = shift_q_map_35;
      end
      6'b100100 : begin
        _zz_shift_q_6_4 = shift_q_map_36;
      end
      6'b100101 : begin
        _zz_shift_q_6_4 = shift_q_map_37;
      end
      6'b100110 : begin
        _zz_shift_q_6_4 = shift_q_map_38;
      end
      default : begin
        _zz_shift_q_6_4 = shift_q_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_7_5)
      6'b000000 : begin
        _zz_shift_i_7_4 = shift_i_map_0;
      end
      6'b000001 : begin
        _zz_shift_i_7_4 = shift_i_map_1;
      end
      6'b000010 : begin
        _zz_shift_i_7_4 = shift_i_map_2;
      end
      6'b000011 : begin
        _zz_shift_i_7_4 = shift_i_map_3;
      end
      6'b000100 : begin
        _zz_shift_i_7_4 = shift_i_map_4;
      end
      6'b000101 : begin
        _zz_shift_i_7_4 = shift_i_map_5;
      end
      6'b000110 : begin
        _zz_shift_i_7_4 = shift_i_map_6;
      end
      6'b000111 : begin
        _zz_shift_i_7_4 = shift_i_map_7;
      end
      6'b001000 : begin
        _zz_shift_i_7_4 = shift_i_map_8;
      end
      6'b001001 : begin
        _zz_shift_i_7_4 = shift_i_map_9;
      end
      6'b001010 : begin
        _zz_shift_i_7_4 = shift_i_map_10;
      end
      6'b001011 : begin
        _zz_shift_i_7_4 = shift_i_map_11;
      end
      6'b001100 : begin
        _zz_shift_i_7_4 = shift_i_map_12;
      end
      6'b001101 : begin
        _zz_shift_i_7_4 = shift_i_map_13;
      end
      6'b001110 : begin
        _zz_shift_i_7_4 = shift_i_map_14;
      end
      6'b001111 : begin
        _zz_shift_i_7_4 = shift_i_map_15;
      end
      6'b010000 : begin
        _zz_shift_i_7_4 = shift_i_map_16;
      end
      6'b010001 : begin
        _zz_shift_i_7_4 = shift_i_map_17;
      end
      6'b010010 : begin
        _zz_shift_i_7_4 = shift_i_map_18;
      end
      6'b010011 : begin
        _zz_shift_i_7_4 = shift_i_map_19;
      end
      6'b010100 : begin
        _zz_shift_i_7_4 = shift_i_map_20;
      end
      6'b010101 : begin
        _zz_shift_i_7_4 = shift_i_map_21;
      end
      6'b010110 : begin
        _zz_shift_i_7_4 = shift_i_map_22;
      end
      6'b010111 : begin
        _zz_shift_i_7_4 = shift_i_map_23;
      end
      6'b011000 : begin
        _zz_shift_i_7_4 = shift_i_map_24;
      end
      6'b011001 : begin
        _zz_shift_i_7_4 = shift_i_map_25;
      end
      6'b011010 : begin
        _zz_shift_i_7_4 = shift_i_map_26;
      end
      6'b011011 : begin
        _zz_shift_i_7_4 = shift_i_map_27;
      end
      6'b011100 : begin
        _zz_shift_i_7_4 = shift_i_map_28;
      end
      6'b011101 : begin
        _zz_shift_i_7_4 = shift_i_map_29;
      end
      6'b011110 : begin
        _zz_shift_i_7_4 = shift_i_map_30;
      end
      6'b011111 : begin
        _zz_shift_i_7_4 = shift_i_map_31;
      end
      6'b100000 : begin
        _zz_shift_i_7_4 = shift_i_map_32;
      end
      6'b100001 : begin
        _zz_shift_i_7_4 = shift_i_map_33;
      end
      6'b100010 : begin
        _zz_shift_i_7_4 = shift_i_map_34;
      end
      6'b100011 : begin
        _zz_shift_i_7_4 = shift_i_map_35;
      end
      6'b100100 : begin
        _zz_shift_i_7_4 = shift_i_map_36;
      end
      6'b100101 : begin
        _zz_shift_i_7_4 = shift_i_map_37;
      end
      6'b100110 : begin
        _zz_shift_i_7_4 = shift_i_map_38;
      end
      default : begin
        _zz_shift_i_7_4 = shift_i_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_7_5)
      6'b000000 : begin
        _zz_shift_q_7_4 = shift_q_map_0;
      end
      6'b000001 : begin
        _zz_shift_q_7_4 = shift_q_map_1;
      end
      6'b000010 : begin
        _zz_shift_q_7_4 = shift_q_map_2;
      end
      6'b000011 : begin
        _zz_shift_q_7_4 = shift_q_map_3;
      end
      6'b000100 : begin
        _zz_shift_q_7_4 = shift_q_map_4;
      end
      6'b000101 : begin
        _zz_shift_q_7_4 = shift_q_map_5;
      end
      6'b000110 : begin
        _zz_shift_q_7_4 = shift_q_map_6;
      end
      6'b000111 : begin
        _zz_shift_q_7_4 = shift_q_map_7;
      end
      6'b001000 : begin
        _zz_shift_q_7_4 = shift_q_map_8;
      end
      6'b001001 : begin
        _zz_shift_q_7_4 = shift_q_map_9;
      end
      6'b001010 : begin
        _zz_shift_q_7_4 = shift_q_map_10;
      end
      6'b001011 : begin
        _zz_shift_q_7_4 = shift_q_map_11;
      end
      6'b001100 : begin
        _zz_shift_q_7_4 = shift_q_map_12;
      end
      6'b001101 : begin
        _zz_shift_q_7_4 = shift_q_map_13;
      end
      6'b001110 : begin
        _zz_shift_q_7_4 = shift_q_map_14;
      end
      6'b001111 : begin
        _zz_shift_q_7_4 = shift_q_map_15;
      end
      6'b010000 : begin
        _zz_shift_q_7_4 = shift_q_map_16;
      end
      6'b010001 : begin
        _zz_shift_q_7_4 = shift_q_map_17;
      end
      6'b010010 : begin
        _zz_shift_q_7_4 = shift_q_map_18;
      end
      6'b010011 : begin
        _zz_shift_q_7_4 = shift_q_map_19;
      end
      6'b010100 : begin
        _zz_shift_q_7_4 = shift_q_map_20;
      end
      6'b010101 : begin
        _zz_shift_q_7_4 = shift_q_map_21;
      end
      6'b010110 : begin
        _zz_shift_q_7_4 = shift_q_map_22;
      end
      6'b010111 : begin
        _zz_shift_q_7_4 = shift_q_map_23;
      end
      6'b011000 : begin
        _zz_shift_q_7_4 = shift_q_map_24;
      end
      6'b011001 : begin
        _zz_shift_q_7_4 = shift_q_map_25;
      end
      6'b011010 : begin
        _zz_shift_q_7_4 = shift_q_map_26;
      end
      6'b011011 : begin
        _zz_shift_q_7_4 = shift_q_map_27;
      end
      6'b011100 : begin
        _zz_shift_q_7_4 = shift_q_map_28;
      end
      6'b011101 : begin
        _zz_shift_q_7_4 = shift_q_map_29;
      end
      6'b011110 : begin
        _zz_shift_q_7_4 = shift_q_map_30;
      end
      6'b011111 : begin
        _zz_shift_q_7_4 = shift_q_map_31;
      end
      6'b100000 : begin
        _zz_shift_q_7_4 = shift_q_map_32;
      end
      6'b100001 : begin
        _zz_shift_q_7_4 = shift_q_map_33;
      end
      6'b100010 : begin
        _zz_shift_q_7_4 = shift_q_map_34;
      end
      6'b100011 : begin
        _zz_shift_q_7_4 = shift_q_map_35;
      end
      6'b100100 : begin
        _zz_shift_q_7_4 = shift_q_map_36;
      end
      6'b100101 : begin
        _zz_shift_q_7_4 = shift_q_map_37;
      end
      6'b100110 : begin
        _zz_shift_q_7_4 = shift_q_map_38;
      end
      default : begin
        _zz_shift_q_7_4 = shift_q_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_0_7)
      6'b000000 : begin
        _zz_shift_i_0_6 = shift_i_map_0;
      end
      6'b000001 : begin
        _zz_shift_i_0_6 = shift_i_map_1;
      end
      6'b000010 : begin
        _zz_shift_i_0_6 = shift_i_map_2;
      end
      6'b000011 : begin
        _zz_shift_i_0_6 = shift_i_map_3;
      end
      6'b000100 : begin
        _zz_shift_i_0_6 = shift_i_map_4;
      end
      6'b000101 : begin
        _zz_shift_i_0_6 = shift_i_map_5;
      end
      6'b000110 : begin
        _zz_shift_i_0_6 = shift_i_map_6;
      end
      6'b000111 : begin
        _zz_shift_i_0_6 = shift_i_map_7;
      end
      6'b001000 : begin
        _zz_shift_i_0_6 = shift_i_map_8;
      end
      6'b001001 : begin
        _zz_shift_i_0_6 = shift_i_map_9;
      end
      6'b001010 : begin
        _zz_shift_i_0_6 = shift_i_map_10;
      end
      6'b001011 : begin
        _zz_shift_i_0_6 = shift_i_map_11;
      end
      6'b001100 : begin
        _zz_shift_i_0_6 = shift_i_map_12;
      end
      6'b001101 : begin
        _zz_shift_i_0_6 = shift_i_map_13;
      end
      6'b001110 : begin
        _zz_shift_i_0_6 = shift_i_map_14;
      end
      6'b001111 : begin
        _zz_shift_i_0_6 = shift_i_map_15;
      end
      6'b010000 : begin
        _zz_shift_i_0_6 = shift_i_map_16;
      end
      6'b010001 : begin
        _zz_shift_i_0_6 = shift_i_map_17;
      end
      6'b010010 : begin
        _zz_shift_i_0_6 = shift_i_map_18;
      end
      6'b010011 : begin
        _zz_shift_i_0_6 = shift_i_map_19;
      end
      6'b010100 : begin
        _zz_shift_i_0_6 = shift_i_map_20;
      end
      6'b010101 : begin
        _zz_shift_i_0_6 = shift_i_map_21;
      end
      6'b010110 : begin
        _zz_shift_i_0_6 = shift_i_map_22;
      end
      6'b010111 : begin
        _zz_shift_i_0_6 = shift_i_map_23;
      end
      6'b011000 : begin
        _zz_shift_i_0_6 = shift_i_map_24;
      end
      6'b011001 : begin
        _zz_shift_i_0_6 = shift_i_map_25;
      end
      6'b011010 : begin
        _zz_shift_i_0_6 = shift_i_map_26;
      end
      6'b011011 : begin
        _zz_shift_i_0_6 = shift_i_map_27;
      end
      6'b011100 : begin
        _zz_shift_i_0_6 = shift_i_map_28;
      end
      6'b011101 : begin
        _zz_shift_i_0_6 = shift_i_map_29;
      end
      6'b011110 : begin
        _zz_shift_i_0_6 = shift_i_map_30;
      end
      6'b011111 : begin
        _zz_shift_i_0_6 = shift_i_map_31;
      end
      6'b100000 : begin
        _zz_shift_i_0_6 = shift_i_map_32;
      end
      6'b100001 : begin
        _zz_shift_i_0_6 = shift_i_map_33;
      end
      6'b100010 : begin
        _zz_shift_i_0_6 = shift_i_map_34;
      end
      6'b100011 : begin
        _zz_shift_i_0_6 = shift_i_map_35;
      end
      6'b100100 : begin
        _zz_shift_i_0_6 = shift_i_map_36;
      end
      6'b100101 : begin
        _zz_shift_i_0_6 = shift_i_map_37;
      end
      6'b100110 : begin
        _zz_shift_i_0_6 = shift_i_map_38;
      end
      default : begin
        _zz_shift_i_0_6 = shift_i_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_0_7)
      6'b000000 : begin
        _zz_shift_q_0_6 = shift_q_map_0;
      end
      6'b000001 : begin
        _zz_shift_q_0_6 = shift_q_map_1;
      end
      6'b000010 : begin
        _zz_shift_q_0_6 = shift_q_map_2;
      end
      6'b000011 : begin
        _zz_shift_q_0_6 = shift_q_map_3;
      end
      6'b000100 : begin
        _zz_shift_q_0_6 = shift_q_map_4;
      end
      6'b000101 : begin
        _zz_shift_q_0_6 = shift_q_map_5;
      end
      6'b000110 : begin
        _zz_shift_q_0_6 = shift_q_map_6;
      end
      6'b000111 : begin
        _zz_shift_q_0_6 = shift_q_map_7;
      end
      6'b001000 : begin
        _zz_shift_q_0_6 = shift_q_map_8;
      end
      6'b001001 : begin
        _zz_shift_q_0_6 = shift_q_map_9;
      end
      6'b001010 : begin
        _zz_shift_q_0_6 = shift_q_map_10;
      end
      6'b001011 : begin
        _zz_shift_q_0_6 = shift_q_map_11;
      end
      6'b001100 : begin
        _zz_shift_q_0_6 = shift_q_map_12;
      end
      6'b001101 : begin
        _zz_shift_q_0_6 = shift_q_map_13;
      end
      6'b001110 : begin
        _zz_shift_q_0_6 = shift_q_map_14;
      end
      6'b001111 : begin
        _zz_shift_q_0_6 = shift_q_map_15;
      end
      6'b010000 : begin
        _zz_shift_q_0_6 = shift_q_map_16;
      end
      6'b010001 : begin
        _zz_shift_q_0_6 = shift_q_map_17;
      end
      6'b010010 : begin
        _zz_shift_q_0_6 = shift_q_map_18;
      end
      6'b010011 : begin
        _zz_shift_q_0_6 = shift_q_map_19;
      end
      6'b010100 : begin
        _zz_shift_q_0_6 = shift_q_map_20;
      end
      6'b010101 : begin
        _zz_shift_q_0_6 = shift_q_map_21;
      end
      6'b010110 : begin
        _zz_shift_q_0_6 = shift_q_map_22;
      end
      6'b010111 : begin
        _zz_shift_q_0_6 = shift_q_map_23;
      end
      6'b011000 : begin
        _zz_shift_q_0_6 = shift_q_map_24;
      end
      6'b011001 : begin
        _zz_shift_q_0_6 = shift_q_map_25;
      end
      6'b011010 : begin
        _zz_shift_q_0_6 = shift_q_map_26;
      end
      6'b011011 : begin
        _zz_shift_q_0_6 = shift_q_map_27;
      end
      6'b011100 : begin
        _zz_shift_q_0_6 = shift_q_map_28;
      end
      6'b011101 : begin
        _zz_shift_q_0_6 = shift_q_map_29;
      end
      6'b011110 : begin
        _zz_shift_q_0_6 = shift_q_map_30;
      end
      6'b011111 : begin
        _zz_shift_q_0_6 = shift_q_map_31;
      end
      6'b100000 : begin
        _zz_shift_q_0_6 = shift_q_map_32;
      end
      6'b100001 : begin
        _zz_shift_q_0_6 = shift_q_map_33;
      end
      6'b100010 : begin
        _zz_shift_q_0_6 = shift_q_map_34;
      end
      6'b100011 : begin
        _zz_shift_q_0_6 = shift_q_map_35;
      end
      6'b100100 : begin
        _zz_shift_q_0_6 = shift_q_map_36;
      end
      6'b100101 : begin
        _zz_shift_q_0_6 = shift_q_map_37;
      end
      6'b100110 : begin
        _zz_shift_q_0_6 = shift_q_map_38;
      end
      default : begin
        _zz_shift_q_0_6 = shift_q_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_1_7)
      6'b000000 : begin
        _zz_shift_i_1_6 = shift_i_map_0;
      end
      6'b000001 : begin
        _zz_shift_i_1_6 = shift_i_map_1;
      end
      6'b000010 : begin
        _zz_shift_i_1_6 = shift_i_map_2;
      end
      6'b000011 : begin
        _zz_shift_i_1_6 = shift_i_map_3;
      end
      6'b000100 : begin
        _zz_shift_i_1_6 = shift_i_map_4;
      end
      6'b000101 : begin
        _zz_shift_i_1_6 = shift_i_map_5;
      end
      6'b000110 : begin
        _zz_shift_i_1_6 = shift_i_map_6;
      end
      6'b000111 : begin
        _zz_shift_i_1_6 = shift_i_map_7;
      end
      6'b001000 : begin
        _zz_shift_i_1_6 = shift_i_map_8;
      end
      6'b001001 : begin
        _zz_shift_i_1_6 = shift_i_map_9;
      end
      6'b001010 : begin
        _zz_shift_i_1_6 = shift_i_map_10;
      end
      6'b001011 : begin
        _zz_shift_i_1_6 = shift_i_map_11;
      end
      6'b001100 : begin
        _zz_shift_i_1_6 = shift_i_map_12;
      end
      6'b001101 : begin
        _zz_shift_i_1_6 = shift_i_map_13;
      end
      6'b001110 : begin
        _zz_shift_i_1_6 = shift_i_map_14;
      end
      6'b001111 : begin
        _zz_shift_i_1_6 = shift_i_map_15;
      end
      6'b010000 : begin
        _zz_shift_i_1_6 = shift_i_map_16;
      end
      6'b010001 : begin
        _zz_shift_i_1_6 = shift_i_map_17;
      end
      6'b010010 : begin
        _zz_shift_i_1_6 = shift_i_map_18;
      end
      6'b010011 : begin
        _zz_shift_i_1_6 = shift_i_map_19;
      end
      6'b010100 : begin
        _zz_shift_i_1_6 = shift_i_map_20;
      end
      6'b010101 : begin
        _zz_shift_i_1_6 = shift_i_map_21;
      end
      6'b010110 : begin
        _zz_shift_i_1_6 = shift_i_map_22;
      end
      6'b010111 : begin
        _zz_shift_i_1_6 = shift_i_map_23;
      end
      6'b011000 : begin
        _zz_shift_i_1_6 = shift_i_map_24;
      end
      6'b011001 : begin
        _zz_shift_i_1_6 = shift_i_map_25;
      end
      6'b011010 : begin
        _zz_shift_i_1_6 = shift_i_map_26;
      end
      6'b011011 : begin
        _zz_shift_i_1_6 = shift_i_map_27;
      end
      6'b011100 : begin
        _zz_shift_i_1_6 = shift_i_map_28;
      end
      6'b011101 : begin
        _zz_shift_i_1_6 = shift_i_map_29;
      end
      6'b011110 : begin
        _zz_shift_i_1_6 = shift_i_map_30;
      end
      6'b011111 : begin
        _zz_shift_i_1_6 = shift_i_map_31;
      end
      6'b100000 : begin
        _zz_shift_i_1_6 = shift_i_map_32;
      end
      6'b100001 : begin
        _zz_shift_i_1_6 = shift_i_map_33;
      end
      6'b100010 : begin
        _zz_shift_i_1_6 = shift_i_map_34;
      end
      6'b100011 : begin
        _zz_shift_i_1_6 = shift_i_map_35;
      end
      6'b100100 : begin
        _zz_shift_i_1_6 = shift_i_map_36;
      end
      6'b100101 : begin
        _zz_shift_i_1_6 = shift_i_map_37;
      end
      6'b100110 : begin
        _zz_shift_i_1_6 = shift_i_map_38;
      end
      default : begin
        _zz_shift_i_1_6 = shift_i_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_1_7)
      6'b000000 : begin
        _zz_shift_q_1_6 = shift_q_map_0;
      end
      6'b000001 : begin
        _zz_shift_q_1_6 = shift_q_map_1;
      end
      6'b000010 : begin
        _zz_shift_q_1_6 = shift_q_map_2;
      end
      6'b000011 : begin
        _zz_shift_q_1_6 = shift_q_map_3;
      end
      6'b000100 : begin
        _zz_shift_q_1_6 = shift_q_map_4;
      end
      6'b000101 : begin
        _zz_shift_q_1_6 = shift_q_map_5;
      end
      6'b000110 : begin
        _zz_shift_q_1_6 = shift_q_map_6;
      end
      6'b000111 : begin
        _zz_shift_q_1_6 = shift_q_map_7;
      end
      6'b001000 : begin
        _zz_shift_q_1_6 = shift_q_map_8;
      end
      6'b001001 : begin
        _zz_shift_q_1_6 = shift_q_map_9;
      end
      6'b001010 : begin
        _zz_shift_q_1_6 = shift_q_map_10;
      end
      6'b001011 : begin
        _zz_shift_q_1_6 = shift_q_map_11;
      end
      6'b001100 : begin
        _zz_shift_q_1_6 = shift_q_map_12;
      end
      6'b001101 : begin
        _zz_shift_q_1_6 = shift_q_map_13;
      end
      6'b001110 : begin
        _zz_shift_q_1_6 = shift_q_map_14;
      end
      6'b001111 : begin
        _zz_shift_q_1_6 = shift_q_map_15;
      end
      6'b010000 : begin
        _zz_shift_q_1_6 = shift_q_map_16;
      end
      6'b010001 : begin
        _zz_shift_q_1_6 = shift_q_map_17;
      end
      6'b010010 : begin
        _zz_shift_q_1_6 = shift_q_map_18;
      end
      6'b010011 : begin
        _zz_shift_q_1_6 = shift_q_map_19;
      end
      6'b010100 : begin
        _zz_shift_q_1_6 = shift_q_map_20;
      end
      6'b010101 : begin
        _zz_shift_q_1_6 = shift_q_map_21;
      end
      6'b010110 : begin
        _zz_shift_q_1_6 = shift_q_map_22;
      end
      6'b010111 : begin
        _zz_shift_q_1_6 = shift_q_map_23;
      end
      6'b011000 : begin
        _zz_shift_q_1_6 = shift_q_map_24;
      end
      6'b011001 : begin
        _zz_shift_q_1_6 = shift_q_map_25;
      end
      6'b011010 : begin
        _zz_shift_q_1_6 = shift_q_map_26;
      end
      6'b011011 : begin
        _zz_shift_q_1_6 = shift_q_map_27;
      end
      6'b011100 : begin
        _zz_shift_q_1_6 = shift_q_map_28;
      end
      6'b011101 : begin
        _zz_shift_q_1_6 = shift_q_map_29;
      end
      6'b011110 : begin
        _zz_shift_q_1_6 = shift_q_map_30;
      end
      6'b011111 : begin
        _zz_shift_q_1_6 = shift_q_map_31;
      end
      6'b100000 : begin
        _zz_shift_q_1_6 = shift_q_map_32;
      end
      6'b100001 : begin
        _zz_shift_q_1_6 = shift_q_map_33;
      end
      6'b100010 : begin
        _zz_shift_q_1_6 = shift_q_map_34;
      end
      6'b100011 : begin
        _zz_shift_q_1_6 = shift_q_map_35;
      end
      6'b100100 : begin
        _zz_shift_q_1_6 = shift_q_map_36;
      end
      6'b100101 : begin
        _zz_shift_q_1_6 = shift_q_map_37;
      end
      6'b100110 : begin
        _zz_shift_q_1_6 = shift_q_map_38;
      end
      default : begin
        _zz_shift_q_1_6 = shift_q_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_2_7)
      6'b000000 : begin
        _zz_shift_i_2_6 = shift_i_map_0;
      end
      6'b000001 : begin
        _zz_shift_i_2_6 = shift_i_map_1;
      end
      6'b000010 : begin
        _zz_shift_i_2_6 = shift_i_map_2;
      end
      6'b000011 : begin
        _zz_shift_i_2_6 = shift_i_map_3;
      end
      6'b000100 : begin
        _zz_shift_i_2_6 = shift_i_map_4;
      end
      6'b000101 : begin
        _zz_shift_i_2_6 = shift_i_map_5;
      end
      6'b000110 : begin
        _zz_shift_i_2_6 = shift_i_map_6;
      end
      6'b000111 : begin
        _zz_shift_i_2_6 = shift_i_map_7;
      end
      6'b001000 : begin
        _zz_shift_i_2_6 = shift_i_map_8;
      end
      6'b001001 : begin
        _zz_shift_i_2_6 = shift_i_map_9;
      end
      6'b001010 : begin
        _zz_shift_i_2_6 = shift_i_map_10;
      end
      6'b001011 : begin
        _zz_shift_i_2_6 = shift_i_map_11;
      end
      6'b001100 : begin
        _zz_shift_i_2_6 = shift_i_map_12;
      end
      6'b001101 : begin
        _zz_shift_i_2_6 = shift_i_map_13;
      end
      6'b001110 : begin
        _zz_shift_i_2_6 = shift_i_map_14;
      end
      6'b001111 : begin
        _zz_shift_i_2_6 = shift_i_map_15;
      end
      6'b010000 : begin
        _zz_shift_i_2_6 = shift_i_map_16;
      end
      6'b010001 : begin
        _zz_shift_i_2_6 = shift_i_map_17;
      end
      6'b010010 : begin
        _zz_shift_i_2_6 = shift_i_map_18;
      end
      6'b010011 : begin
        _zz_shift_i_2_6 = shift_i_map_19;
      end
      6'b010100 : begin
        _zz_shift_i_2_6 = shift_i_map_20;
      end
      6'b010101 : begin
        _zz_shift_i_2_6 = shift_i_map_21;
      end
      6'b010110 : begin
        _zz_shift_i_2_6 = shift_i_map_22;
      end
      6'b010111 : begin
        _zz_shift_i_2_6 = shift_i_map_23;
      end
      6'b011000 : begin
        _zz_shift_i_2_6 = shift_i_map_24;
      end
      6'b011001 : begin
        _zz_shift_i_2_6 = shift_i_map_25;
      end
      6'b011010 : begin
        _zz_shift_i_2_6 = shift_i_map_26;
      end
      6'b011011 : begin
        _zz_shift_i_2_6 = shift_i_map_27;
      end
      6'b011100 : begin
        _zz_shift_i_2_6 = shift_i_map_28;
      end
      6'b011101 : begin
        _zz_shift_i_2_6 = shift_i_map_29;
      end
      6'b011110 : begin
        _zz_shift_i_2_6 = shift_i_map_30;
      end
      6'b011111 : begin
        _zz_shift_i_2_6 = shift_i_map_31;
      end
      6'b100000 : begin
        _zz_shift_i_2_6 = shift_i_map_32;
      end
      6'b100001 : begin
        _zz_shift_i_2_6 = shift_i_map_33;
      end
      6'b100010 : begin
        _zz_shift_i_2_6 = shift_i_map_34;
      end
      6'b100011 : begin
        _zz_shift_i_2_6 = shift_i_map_35;
      end
      6'b100100 : begin
        _zz_shift_i_2_6 = shift_i_map_36;
      end
      6'b100101 : begin
        _zz_shift_i_2_6 = shift_i_map_37;
      end
      6'b100110 : begin
        _zz_shift_i_2_6 = shift_i_map_38;
      end
      default : begin
        _zz_shift_i_2_6 = shift_i_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_2_7)
      6'b000000 : begin
        _zz_shift_q_2_6 = shift_q_map_0;
      end
      6'b000001 : begin
        _zz_shift_q_2_6 = shift_q_map_1;
      end
      6'b000010 : begin
        _zz_shift_q_2_6 = shift_q_map_2;
      end
      6'b000011 : begin
        _zz_shift_q_2_6 = shift_q_map_3;
      end
      6'b000100 : begin
        _zz_shift_q_2_6 = shift_q_map_4;
      end
      6'b000101 : begin
        _zz_shift_q_2_6 = shift_q_map_5;
      end
      6'b000110 : begin
        _zz_shift_q_2_6 = shift_q_map_6;
      end
      6'b000111 : begin
        _zz_shift_q_2_6 = shift_q_map_7;
      end
      6'b001000 : begin
        _zz_shift_q_2_6 = shift_q_map_8;
      end
      6'b001001 : begin
        _zz_shift_q_2_6 = shift_q_map_9;
      end
      6'b001010 : begin
        _zz_shift_q_2_6 = shift_q_map_10;
      end
      6'b001011 : begin
        _zz_shift_q_2_6 = shift_q_map_11;
      end
      6'b001100 : begin
        _zz_shift_q_2_6 = shift_q_map_12;
      end
      6'b001101 : begin
        _zz_shift_q_2_6 = shift_q_map_13;
      end
      6'b001110 : begin
        _zz_shift_q_2_6 = shift_q_map_14;
      end
      6'b001111 : begin
        _zz_shift_q_2_6 = shift_q_map_15;
      end
      6'b010000 : begin
        _zz_shift_q_2_6 = shift_q_map_16;
      end
      6'b010001 : begin
        _zz_shift_q_2_6 = shift_q_map_17;
      end
      6'b010010 : begin
        _zz_shift_q_2_6 = shift_q_map_18;
      end
      6'b010011 : begin
        _zz_shift_q_2_6 = shift_q_map_19;
      end
      6'b010100 : begin
        _zz_shift_q_2_6 = shift_q_map_20;
      end
      6'b010101 : begin
        _zz_shift_q_2_6 = shift_q_map_21;
      end
      6'b010110 : begin
        _zz_shift_q_2_6 = shift_q_map_22;
      end
      6'b010111 : begin
        _zz_shift_q_2_6 = shift_q_map_23;
      end
      6'b011000 : begin
        _zz_shift_q_2_6 = shift_q_map_24;
      end
      6'b011001 : begin
        _zz_shift_q_2_6 = shift_q_map_25;
      end
      6'b011010 : begin
        _zz_shift_q_2_6 = shift_q_map_26;
      end
      6'b011011 : begin
        _zz_shift_q_2_6 = shift_q_map_27;
      end
      6'b011100 : begin
        _zz_shift_q_2_6 = shift_q_map_28;
      end
      6'b011101 : begin
        _zz_shift_q_2_6 = shift_q_map_29;
      end
      6'b011110 : begin
        _zz_shift_q_2_6 = shift_q_map_30;
      end
      6'b011111 : begin
        _zz_shift_q_2_6 = shift_q_map_31;
      end
      6'b100000 : begin
        _zz_shift_q_2_6 = shift_q_map_32;
      end
      6'b100001 : begin
        _zz_shift_q_2_6 = shift_q_map_33;
      end
      6'b100010 : begin
        _zz_shift_q_2_6 = shift_q_map_34;
      end
      6'b100011 : begin
        _zz_shift_q_2_6 = shift_q_map_35;
      end
      6'b100100 : begin
        _zz_shift_q_2_6 = shift_q_map_36;
      end
      6'b100101 : begin
        _zz_shift_q_2_6 = shift_q_map_37;
      end
      6'b100110 : begin
        _zz_shift_q_2_6 = shift_q_map_38;
      end
      default : begin
        _zz_shift_q_2_6 = shift_q_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_3_7)
      6'b000000 : begin
        _zz_shift_i_3_6 = shift_i_map_0;
      end
      6'b000001 : begin
        _zz_shift_i_3_6 = shift_i_map_1;
      end
      6'b000010 : begin
        _zz_shift_i_3_6 = shift_i_map_2;
      end
      6'b000011 : begin
        _zz_shift_i_3_6 = shift_i_map_3;
      end
      6'b000100 : begin
        _zz_shift_i_3_6 = shift_i_map_4;
      end
      6'b000101 : begin
        _zz_shift_i_3_6 = shift_i_map_5;
      end
      6'b000110 : begin
        _zz_shift_i_3_6 = shift_i_map_6;
      end
      6'b000111 : begin
        _zz_shift_i_3_6 = shift_i_map_7;
      end
      6'b001000 : begin
        _zz_shift_i_3_6 = shift_i_map_8;
      end
      6'b001001 : begin
        _zz_shift_i_3_6 = shift_i_map_9;
      end
      6'b001010 : begin
        _zz_shift_i_3_6 = shift_i_map_10;
      end
      6'b001011 : begin
        _zz_shift_i_3_6 = shift_i_map_11;
      end
      6'b001100 : begin
        _zz_shift_i_3_6 = shift_i_map_12;
      end
      6'b001101 : begin
        _zz_shift_i_3_6 = shift_i_map_13;
      end
      6'b001110 : begin
        _zz_shift_i_3_6 = shift_i_map_14;
      end
      6'b001111 : begin
        _zz_shift_i_3_6 = shift_i_map_15;
      end
      6'b010000 : begin
        _zz_shift_i_3_6 = shift_i_map_16;
      end
      6'b010001 : begin
        _zz_shift_i_3_6 = shift_i_map_17;
      end
      6'b010010 : begin
        _zz_shift_i_3_6 = shift_i_map_18;
      end
      6'b010011 : begin
        _zz_shift_i_3_6 = shift_i_map_19;
      end
      6'b010100 : begin
        _zz_shift_i_3_6 = shift_i_map_20;
      end
      6'b010101 : begin
        _zz_shift_i_3_6 = shift_i_map_21;
      end
      6'b010110 : begin
        _zz_shift_i_3_6 = shift_i_map_22;
      end
      6'b010111 : begin
        _zz_shift_i_3_6 = shift_i_map_23;
      end
      6'b011000 : begin
        _zz_shift_i_3_6 = shift_i_map_24;
      end
      6'b011001 : begin
        _zz_shift_i_3_6 = shift_i_map_25;
      end
      6'b011010 : begin
        _zz_shift_i_3_6 = shift_i_map_26;
      end
      6'b011011 : begin
        _zz_shift_i_3_6 = shift_i_map_27;
      end
      6'b011100 : begin
        _zz_shift_i_3_6 = shift_i_map_28;
      end
      6'b011101 : begin
        _zz_shift_i_3_6 = shift_i_map_29;
      end
      6'b011110 : begin
        _zz_shift_i_3_6 = shift_i_map_30;
      end
      6'b011111 : begin
        _zz_shift_i_3_6 = shift_i_map_31;
      end
      6'b100000 : begin
        _zz_shift_i_3_6 = shift_i_map_32;
      end
      6'b100001 : begin
        _zz_shift_i_3_6 = shift_i_map_33;
      end
      6'b100010 : begin
        _zz_shift_i_3_6 = shift_i_map_34;
      end
      6'b100011 : begin
        _zz_shift_i_3_6 = shift_i_map_35;
      end
      6'b100100 : begin
        _zz_shift_i_3_6 = shift_i_map_36;
      end
      6'b100101 : begin
        _zz_shift_i_3_6 = shift_i_map_37;
      end
      6'b100110 : begin
        _zz_shift_i_3_6 = shift_i_map_38;
      end
      default : begin
        _zz_shift_i_3_6 = shift_i_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_3_7)
      6'b000000 : begin
        _zz_shift_q_3_6 = shift_q_map_0;
      end
      6'b000001 : begin
        _zz_shift_q_3_6 = shift_q_map_1;
      end
      6'b000010 : begin
        _zz_shift_q_3_6 = shift_q_map_2;
      end
      6'b000011 : begin
        _zz_shift_q_3_6 = shift_q_map_3;
      end
      6'b000100 : begin
        _zz_shift_q_3_6 = shift_q_map_4;
      end
      6'b000101 : begin
        _zz_shift_q_3_6 = shift_q_map_5;
      end
      6'b000110 : begin
        _zz_shift_q_3_6 = shift_q_map_6;
      end
      6'b000111 : begin
        _zz_shift_q_3_6 = shift_q_map_7;
      end
      6'b001000 : begin
        _zz_shift_q_3_6 = shift_q_map_8;
      end
      6'b001001 : begin
        _zz_shift_q_3_6 = shift_q_map_9;
      end
      6'b001010 : begin
        _zz_shift_q_3_6 = shift_q_map_10;
      end
      6'b001011 : begin
        _zz_shift_q_3_6 = shift_q_map_11;
      end
      6'b001100 : begin
        _zz_shift_q_3_6 = shift_q_map_12;
      end
      6'b001101 : begin
        _zz_shift_q_3_6 = shift_q_map_13;
      end
      6'b001110 : begin
        _zz_shift_q_3_6 = shift_q_map_14;
      end
      6'b001111 : begin
        _zz_shift_q_3_6 = shift_q_map_15;
      end
      6'b010000 : begin
        _zz_shift_q_3_6 = shift_q_map_16;
      end
      6'b010001 : begin
        _zz_shift_q_3_6 = shift_q_map_17;
      end
      6'b010010 : begin
        _zz_shift_q_3_6 = shift_q_map_18;
      end
      6'b010011 : begin
        _zz_shift_q_3_6 = shift_q_map_19;
      end
      6'b010100 : begin
        _zz_shift_q_3_6 = shift_q_map_20;
      end
      6'b010101 : begin
        _zz_shift_q_3_6 = shift_q_map_21;
      end
      6'b010110 : begin
        _zz_shift_q_3_6 = shift_q_map_22;
      end
      6'b010111 : begin
        _zz_shift_q_3_6 = shift_q_map_23;
      end
      6'b011000 : begin
        _zz_shift_q_3_6 = shift_q_map_24;
      end
      6'b011001 : begin
        _zz_shift_q_3_6 = shift_q_map_25;
      end
      6'b011010 : begin
        _zz_shift_q_3_6 = shift_q_map_26;
      end
      6'b011011 : begin
        _zz_shift_q_3_6 = shift_q_map_27;
      end
      6'b011100 : begin
        _zz_shift_q_3_6 = shift_q_map_28;
      end
      6'b011101 : begin
        _zz_shift_q_3_6 = shift_q_map_29;
      end
      6'b011110 : begin
        _zz_shift_q_3_6 = shift_q_map_30;
      end
      6'b011111 : begin
        _zz_shift_q_3_6 = shift_q_map_31;
      end
      6'b100000 : begin
        _zz_shift_q_3_6 = shift_q_map_32;
      end
      6'b100001 : begin
        _zz_shift_q_3_6 = shift_q_map_33;
      end
      6'b100010 : begin
        _zz_shift_q_3_6 = shift_q_map_34;
      end
      6'b100011 : begin
        _zz_shift_q_3_6 = shift_q_map_35;
      end
      6'b100100 : begin
        _zz_shift_q_3_6 = shift_q_map_36;
      end
      6'b100101 : begin
        _zz_shift_q_3_6 = shift_q_map_37;
      end
      6'b100110 : begin
        _zz_shift_q_3_6 = shift_q_map_38;
      end
      default : begin
        _zz_shift_q_3_6 = shift_q_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_4_7)
      6'b000000 : begin
        _zz_shift_i_4_6 = shift_i_map_0;
      end
      6'b000001 : begin
        _zz_shift_i_4_6 = shift_i_map_1;
      end
      6'b000010 : begin
        _zz_shift_i_4_6 = shift_i_map_2;
      end
      6'b000011 : begin
        _zz_shift_i_4_6 = shift_i_map_3;
      end
      6'b000100 : begin
        _zz_shift_i_4_6 = shift_i_map_4;
      end
      6'b000101 : begin
        _zz_shift_i_4_6 = shift_i_map_5;
      end
      6'b000110 : begin
        _zz_shift_i_4_6 = shift_i_map_6;
      end
      6'b000111 : begin
        _zz_shift_i_4_6 = shift_i_map_7;
      end
      6'b001000 : begin
        _zz_shift_i_4_6 = shift_i_map_8;
      end
      6'b001001 : begin
        _zz_shift_i_4_6 = shift_i_map_9;
      end
      6'b001010 : begin
        _zz_shift_i_4_6 = shift_i_map_10;
      end
      6'b001011 : begin
        _zz_shift_i_4_6 = shift_i_map_11;
      end
      6'b001100 : begin
        _zz_shift_i_4_6 = shift_i_map_12;
      end
      6'b001101 : begin
        _zz_shift_i_4_6 = shift_i_map_13;
      end
      6'b001110 : begin
        _zz_shift_i_4_6 = shift_i_map_14;
      end
      6'b001111 : begin
        _zz_shift_i_4_6 = shift_i_map_15;
      end
      6'b010000 : begin
        _zz_shift_i_4_6 = shift_i_map_16;
      end
      6'b010001 : begin
        _zz_shift_i_4_6 = shift_i_map_17;
      end
      6'b010010 : begin
        _zz_shift_i_4_6 = shift_i_map_18;
      end
      6'b010011 : begin
        _zz_shift_i_4_6 = shift_i_map_19;
      end
      6'b010100 : begin
        _zz_shift_i_4_6 = shift_i_map_20;
      end
      6'b010101 : begin
        _zz_shift_i_4_6 = shift_i_map_21;
      end
      6'b010110 : begin
        _zz_shift_i_4_6 = shift_i_map_22;
      end
      6'b010111 : begin
        _zz_shift_i_4_6 = shift_i_map_23;
      end
      6'b011000 : begin
        _zz_shift_i_4_6 = shift_i_map_24;
      end
      6'b011001 : begin
        _zz_shift_i_4_6 = shift_i_map_25;
      end
      6'b011010 : begin
        _zz_shift_i_4_6 = shift_i_map_26;
      end
      6'b011011 : begin
        _zz_shift_i_4_6 = shift_i_map_27;
      end
      6'b011100 : begin
        _zz_shift_i_4_6 = shift_i_map_28;
      end
      6'b011101 : begin
        _zz_shift_i_4_6 = shift_i_map_29;
      end
      6'b011110 : begin
        _zz_shift_i_4_6 = shift_i_map_30;
      end
      6'b011111 : begin
        _zz_shift_i_4_6 = shift_i_map_31;
      end
      6'b100000 : begin
        _zz_shift_i_4_6 = shift_i_map_32;
      end
      6'b100001 : begin
        _zz_shift_i_4_6 = shift_i_map_33;
      end
      6'b100010 : begin
        _zz_shift_i_4_6 = shift_i_map_34;
      end
      6'b100011 : begin
        _zz_shift_i_4_6 = shift_i_map_35;
      end
      6'b100100 : begin
        _zz_shift_i_4_6 = shift_i_map_36;
      end
      6'b100101 : begin
        _zz_shift_i_4_6 = shift_i_map_37;
      end
      6'b100110 : begin
        _zz_shift_i_4_6 = shift_i_map_38;
      end
      default : begin
        _zz_shift_i_4_6 = shift_i_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_4_7)
      6'b000000 : begin
        _zz_shift_q_4_6 = shift_q_map_0;
      end
      6'b000001 : begin
        _zz_shift_q_4_6 = shift_q_map_1;
      end
      6'b000010 : begin
        _zz_shift_q_4_6 = shift_q_map_2;
      end
      6'b000011 : begin
        _zz_shift_q_4_6 = shift_q_map_3;
      end
      6'b000100 : begin
        _zz_shift_q_4_6 = shift_q_map_4;
      end
      6'b000101 : begin
        _zz_shift_q_4_6 = shift_q_map_5;
      end
      6'b000110 : begin
        _zz_shift_q_4_6 = shift_q_map_6;
      end
      6'b000111 : begin
        _zz_shift_q_4_6 = shift_q_map_7;
      end
      6'b001000 : begin
        _zz_shift_q_4_6 = shift_q_map_8;
      end
      6'b001001 : begin
        _zz_shift_q_4_6 = shift_q_map_9;
      end
      6'b001010 : begin
        _zz_shift_q_4_6 = shift_q_map_10;
      end
      6'b001011 : begin
        _zz_shift_q_4_6 = shift_q_map_11;
      end
      6'b001100 : begin
        _zz_shift_q_4_6 = shift_q_map_12;
      end
      6'b001101 : begin
        _zz_shift_q_4_6 = shift_q_map_13;
      end
      6'b001110 : begin
        _zz_shift_q_4_6 = shift_q_map_14;
      end
      6'b001111 : begin
        _zz_shift_q_4_6 = shift_q_map_15;
      end
      6'b010000 : begin
        _zz_shift_q_4_6 = shift_q_map_16;
      end
      6'b010001 : begin
        _zz_shift_q_4_6 = shift_q_map_17;
      end
      6'b010010 : begin
        _zz_shift_q_4_6 = shift_q_map_18;
      end
      6'b010011 : begin
        _zz_shift_q_4_6 = shift_q_map_19;
      end
      6'b010100 : begin
        _zz_shift_q_4_6 = shift_q_map_20;
      end
      6'b010101 : begin
        _zz_shift_q_4_6 = shift_q_map_21;
      end
      6'b010110 : begin
        _zz_shift_q_4_6 = shift_q_map_22;
      end
      6'b010111 : begin
        _zz_shift_q_4_6 = shift_q_map_23;
      end
      6'b011000 : begin
        _zz_shift_q_4_6 = shift_q_map_24;
      end
      6'b011001 : begin
        _zz_shift_q_4_6 = shift_q_map_25;
      end
      6'b011010 : begin
        _zz_shift_q_4_6 = shift_q_map_26;
      end
      6'b011011 : begin
        _zz_shift_q_4_6 = shift_q_map_27;
      end
      6'b011100 : begin
        _zz_shift_q_4_6 = shift_q_map_28;
      end
      6'b011101 : begin
        _zz_shift_q_4_6 = shift_q_map_29;
      end
      6'b011110 : begin
        _zz_shift_q_4_6 = shift_q_map_30;
      end
      6'b011111 : begin
        _zz_shift_q_4_6 = shift_q_map_31;
      end
      6'b100000 : begin
        _zz_shift_q_4_6 = shift_q_map_32;
      end
      6'b100001 : begin
        _zz_shift_q_4_6 = shift_q_map_33;
      end
      6'b100010 : begin
        _zz_shift_q_4_6 = shift_q_map_34;
      end
      6'b100011 : begin
        _zz_shift_q_4_6 = shift_q_map_35;
      end
      6'b100100 : begin
        _zz_shift_q_4_6 = shift_q_map_36;
      end
      6'b100101 : begin
        _zz_shift_q_4_6 = shift_q_map_37;
      end
      6'b100110 : begin
        _zz_shift_q_4_6 = shift_q_map_38;
      end
      default : begin
        _zz_shift_q_4_6 = shift_q_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_5_7)
      6'b000000 : begin
        _zz_shift_i_5_6 = shift_i_map_0;
      end
      6'b000001 : begin
        _zz_shift_i_5_6 = shift_i_map_1;
      end
      6'b000010 : begin
        _zz_shift_i_5_6 = shift_i_map_2;
      end
      6'b000011 : begin
        _zz_shift_i_5_6 = shift_i_map_3;
      end
      6'b000100 : begin
        _zz_shift_i_5_6 = shift_i_map_4;
      end
      6'b000101 : begin
        _zz_shift_i_5_6 = shift_i_map_5;
      end
      6'b000110 : begin
        _zz_shift_i_5_6 = shift_i_map_6;
      end
      6'b000111 : begin
        _zz_shift_i_5_6 = shift_i_map_7;
      end
      6'b001000 : begin
        _zz_shift_i_5_6 = shift_i_map_8;
      end
      6'b001001 : begin
        _zz_shift_i_5_6 = shift_i_map_9;
      end
      6'b001010 : begin
        _zz_shift_i_5_6 = shift_i_map_10;
      end
      6'b001011 : begin
        _zz_shift_i_5_6 = shift_i_map_11;
      end
      6'b001100 : begin
        _zz_shift_i_5_6 = shift_i_map_12;
      end
      6'b001101 : begin
        _zz_shift_i_5_6 = shift_i_map_13;
      end
      6'b001110 : begin
        _zz_shift_i_5_6 = shift_i_map_14;
      end
      6'b001111 : begin
        _zz_shift_i_5_6 = shift_i_map_15;
      end
      6'b010000 : begin
        _zz_shift_i_5_6 = shift_i_map_16;
      end
      6'b010001 : begin
        _zz_shift_i_5_6 = shift_i_map_17;
      end
      6'b010010 : begin
        _zz_shift_i_5_6 = shift_i_map_18;
      end
      6'b010011 : begin
        _zz_shift_i_5_6 = shift_i_map_19;
      end
      6'b010100 : begin
        _zz_shift_i_5_6 = shift_i_map_20;
      end
      6'b010101 : begin
        _zz_shift_i_5_6 = shift_i_map_21;
      end
      6'b010110 : begin
        _zz_shift_i_5_6 = shift_i_map_22;
      end
      6'b010111 : begin
        _zz_shift_i_5_6 = shift_i_map_23;
      end
      6'b011000 : begin
        _zz_shift_i_5_6 = shift_i_map_24;
      end
      6'b011001 : begin
        _zz_shift_i_5_6 = shift_i_map_25;
      end
      6'b011010 : begin
        _zz_shift_i_5_6 = shift_i_map_26;
      end
      6'b011011 : begin
        _zz_shift_i_5_6 = shift_i_map_27;
      end
      6'b011100 : begin
        _zz_shift_i_5_6 = shift_i_map_28;
      end
      6'b011101 : begin
        _zz_shift_i_5_6 = shift_i_map_29;
      end
      6'b011110 : begin
        _zz_shift_i_5_6 = shift_i_map_30;
      end
      6'b011111 : begin
        _zz_shift_i_5_6 = shift_i_map_31;
      end
      6'b100000 : begin
        _zz_shift_i_5_6 = shift_i_map_32;
      end
      6'b100001 : begin
        _zz_shift_i_5_6 = shift_i_map_33;
      end
      6'b100010 : begin
        _zz_shift_i_5_6 = shift_i_map_34;
      end
      6'b100011 : begin
        _zz_shift_i_5_6 = shift_i_map_35;
      end
      6'b100100 : begin
        _zz_shift_i_5_6 = shift_i_map_36;
      end
      6'b100101 : begin
        _zz_shift_i_5_6 = shift_i_map_37;
      end
      6'b100110 : begin
        _zz_shift_i_5_6 = shift_i_map_38;
      end
      default : begin
        _zz_shift_i_5_6 = shift_i_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_5_7)
      6'b000000 : begin
        _zz_shift_q_5_6 = shift_q_map_0;
      end
      6'b000001 : begin
        _zz_shift_q_5_6 = shift_q_map_1;
      end
      6'b000010 : begin
        _zz_shift_q_5_6 = shift_q_map_2;
      end
      6'b000011 : begin
        _zz_shift_q_5_6 = shift_q_map_3;
      end
      6'b000100 : begin
        _zz_shift_q_5_6 = shift_q_map_4;
      end
      6'b000101 : begin
        _zz_shift_q_5_6 = shift_q_map_5;
      end
      6'b000110 : begin
        _zz_shift_q_5_6 = shift_q_map_6;
      end
      6'b000111 : begin
        _zz_shift_q_5_6 = shift_q_map_7;
      end
      6'b001000 : begin
        _zz_shift_q_5_6 = shift_q_map_8;
      end
      6'b001001 : begin
        _zz_shift_q_5_6 = shift_q_map_9;
      end
      6'b001010 : begin
        _zz_shift_q_5_6 = shift_q_map_10;
      end
      6'b001011 : begin
        _zz_shift_q_5_6 = shift_q_map_11;
      end
      6'b001100 : begin
        _zz_shift_q_5_6 = shift_q_map_12;
      end
      6'b001101 : begin
        _zz_shift_q_5_6 = shift_q_map_13;
      end
      6'b001110 : begin
        _zz_shift_q_5_6 = shift_q_map_14;
      end
      6'b001111 : begin
        _zz_shift_q_5_6 = shift_q_map_15;
      end
      6'b010000 : begin
        _zz_shift_q_5_6 = shift_q_map_16;
      end
      6'b010001 : begin
        _zz_shift_q_5_6 = shift_q_map_17;
      end
      6'b010010 : begin
        _zz_shift_q_5_6 = shift_q_map_18;
      end
      6'b010011 : begin
        _zz_shift_q_5_6 = shift_q_map_19;
      end
      6'b010100 : begin
        _zz_shift_q_5_6 = shift_q_map_20;
      end
      6'b010101 : begin
        _zz_shift_q_5_6 = shift_q_map_21;
      end
      6'b010110 : begin
        _zz_shift_q_5_6 = shift_q_map_22;
      end
      6'b010111 : begin
        _zz_shift_q_5_6 = shift_q_map_23;
      end
      6'b011000 : begin
        _zz_shift_q_5_6 = shift_q_map_24;
      end
      6'b011001 : begin
        _zz_shift_q_5_6 = shift_q_map_25;
      end
      6'b011010 : begin
        _zz_shift_q_5_6 = shift_q_map_26;
      end
      6'b011011 : begin
        _zz_shift_q_5_6 = shift_q_map_27;
      end
      6'b011100 : begin
        _zz_shift_q_5_6 = shift_q_map_28;
      end
      6'b011101 : begin
        _zz_shift_q_5_6 = shift_q_map_29;
      end
      6'b011110 : begin
        _zz_shift_q_5_6 = shift_q_map_30;
      end
      6'b011111 : begin
        _zz_shift_q_5_6 = shift_q_map_31;
      end
      6'b100000 : begin
        _zz_shift_q_5_6 = shift_q_map_32;
      end
      6'b100001 : begin
        _zz_shift_q_5_6 = shift_q_map_33;
      end
      6'b100010 : begin
        _zz_shift_q_5_6 = shift_q_map_34;
      end
      6'b100011 : begin
        _zz_shift_q_5_6 = shift_q_map_35;
      end
      6'b100100 : begin
        _zz_shift_q_5_6 = shift_q_map_36;
      end
      6'b100101 : begin
        _zz_shift_q_5_6 = shift_q_map_37;
      end
      6'b100110 : begin
        _zz_shift_q_5_6 = shift_q_map_38;
      end
      default : begin
        _zz_shift_q_5_6 = shift_q_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_6_7)
      6'b000000 : begin
        _zz_shift_i_6_6 = shift_i_map_0;
      end
      6'b000001 : begin
        _zz_shift_i_6_6 = shift_i_map_1;
      end
      6'b000010 : begin
        _zz_shift_i_6_6 = shift_i_map_2;
      end
      6'b000011 : begin
        _zz_shift_i_6_6 = shift_i_map_3;
      end
      6'b000100 : begin
        _zz_shift_i_6_6 = shift_i_map_4;
      end
      6'b000101 : begin
        _zz_shift_i_6_6 = shift_i_map_5;
      end
      6'b000110 : begin
        _zz_shift_i_6_6 = shift_i_map_6;
      end
      6'b000111 : begin
        _zz_shift_i_6_6 = shift_i_map_7;
      end
      6'b001000 : begin
        _zz_shift_i_6_6 = shift_i_map_8;
      end
      6'b001001 : begin
        _zz_shift_i_6_6 = shift_i_map_9;
      end
      6'b001010 : begin
        _zz_shift_i_6_6 = shift_i_map_10;
      end
      6'b001011 : begin
        _zz_shift_i_6_6 = shift_i_map_11;
      end
      6'b001100 : begin
        _zz_shift_i_6_6 = shift_i_map_12;
      end
      6'b001101 : begin
        _zz_shift_i_6_6 = shift_i_map_13;
      end
      6'b001110 : begin
        _zz_shift_i_6_6 = shift_i_map_14;
      end
      6'b001111 : begin
        _zz_shift_i_6_6 = shift_i_map_15;
      end
      6'b010000 : begin
        _zz_shift_i_6_6 = shift_i_map_16;
      end
      6'b010001 : begin
        _zz_shift_i_6_6 = shift_i_map_17;
      end
      6'b010010 : begin
        _zz_shift_i_6_6 = shift_i_map_18;
      end
      6'b010011 : begin
        _zz_shift_i_6_6 = shift_i_map_19;
      end
      6'b010100 : begin
        _zz_shift_i_6_6 = shift_i_map_20;
      end
      6'b010101 : begin
        _zz_shift_i_6_6 = shift_i_map_21;
      end
      6'b010110 : begin
        _zz_shift_i_6_6 = shift_i_map_22;
      end
      6'b010111 : begin
        _zz_shift_i_6_6 = shift_i_map_23;
      end
      6'b011000 : begin
        _zz_shift_i_6_6 = shift_i_map_24;
      end
      6'b011001 : begin
        _zz_shift_i_6_6 = shift_i_map_25;
      end
      6'b011010 : begin
        _zz_shift_i_6_6 = shift_i_map_26;
      end
      6'b011011 : begin
        _zz_shift_i_6_6 = shift_i_map_27;
      end
      6'b011100 : begin
        _zz_shift_i_6_6 = shift_i_map_28;
      end
      6'b011101 : begin
        _zz_shift_i_6_6 = shift_i_map_29;
      end
      6'b011110 : begin
        _zz_shift_i_6_6 = shift_i_map_30;
      end
      6'b011111 : begin
        _zz_shift_i_6_6 = shift_i_map_31;
      end
      6'b100000 : begin
        _zz_shift_i_6_6 = shift_i_map_32;
      end
      6'b100001 : begin
        _zz_shift_i_6_6 = shift_i_map_33;
      end
      6'b100010 : begin
        _zz_shift_i_6_6 = shift_i_map_34;
      end
      6'b100011 : begin
        _zz_shift_i_6_6 = shift_i_map_35;
      end
      6'b100100 : begin
        _zz_shift_i_6_6 = shift_i_map_36;
      end
      6'b100101 : begin
        _zz_shift_i_6_6 = shift_i_map_37;
      end
      6'b100110 : begin
        _zz_shift_i_6_6 = shift_i_map_38;
      end
      default : begin
        _zz_shift_i_6_6 = shift_i_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_6_7)
      6'b000000 : begin
        _zz_shift_q_6_6 = shift_q_map_0;
      end
      6'b000001 : begin
        _zz_shift_q_6_6 = shift_q_map_1;
      end
      6'b000010 : begin
        _zz_shift_q_6_6 = shift_q_map_2;
      end
      6'b000011 : begin
        _zz_shift_q_6_6 = shift_q_map_3;
      end
      6'b000100 : begin
        _zz_shift_q_6_6 = shift_q_map_4;
      end
      6'b000101 : begin
        _zz_shift_q_6_6 = shift_q_map_5;
      end
      6'b000110 : begin
        _zz_shift_q_6_6 = shift_q_map_6;
      end
      6'b000111 : begin
        _zz_shift_q_6_6 = shift_q_map_7;
      end
      6'b001000 : begin
        _zz_shift_q_6_6 = shift_q_map_8;
      end
      6'b001001 : begin
        _zz_shift_q_6_6 = shift_q_map_9;
      end
      6'b001010 : begin
        _zz_shift_q_6_6 = shift_q_map_10;
      end
      6'b001011 : begin
        _zz_shift_q_6_6 = shift_q_map_11;
      end
      6'b001100 : begin
        _zz_shift_q_6_6 = shift_q_map_12;
      end
      6'b001101 : begin
        _zz_shift_q_6_6 = shift_q_map_13;
      end
      6'b001110 : begin
        _zz_shift_q_6_6 = shift_q_map_14;
      end
      6'b001111 : begin
        _zz_shift_q_6_6 = shift_q_map_15;
      end
      6'b010000 : begin
        _zz_shift_q_6_6 = shift_q_map_16;
      end
      6'b010001 : begin
        _zz_shift_q_6_6 = shift_q_map_17;
      end
      6'b010010 : begin
        _zz_shift_q_6_6 = shift_q_map_18;
      end
      6'b010011 : begin
        _zz_shift_q_6_6 = shift_q_map_19;
      end
      6'b010100 : begin
        _zz_shift_q_6_6 = shift_q_map_20;
      end
      6'b010101 : begin
        _zz_shift_q_6_6 = shift_q_map_21;
      end
      6'b010110 : begin
        _zz_shift_q_6_6 = shift_q_map_22;
      end
      6'b010111 : begin
        _zz_shift_q_6_6 = shift_q_map_23;
      end
      6'b011000 : begin
        _zz_shift_q_6_6 = shift_q_map_24;
      end
      6'b011001 : begin
        _zz_shift_q_6_6 = shift_q_map_25;
      end
      6'b011010 : begin
        _zz_shift_q_6_6 = shift_q_map_26;
      end
      6'b011011 : begin
        _zz_shift_q_6_6 = shift_q_map_27;
      end
      6'b011100 : begin
        _zz_shift_q_6_6 = shift_q_map_28;
      end
      6'b011101 : begin
        _zz_shift_q_6_6 = shift_q_map_29;
      end
      6'b011110 : begin
        _zz_shift_q_6_6 = shift_q_map_30;
      end
      6'b011111 : begin
        _zz_shift_q_6_6 = shift_q_map_31;
      end
      6'b100000 : begin
        _zz_shift_q_6_6 = shift_q_map_32;
      end
      6'b100001 : begin
        _zz_shift_q_6_6 = shift_q_map_33;
      end
      6'b100010 : begin
        _zz_shift_q_6_6 = shift_q_map_34;
      end
      6'b100011 : begin
        _zz_shift_q_6_6 = shift_q_map_35;
      end
      6'b100100 : begin
        _zz_shift_q_6_6 = shift_q_map_36;
      end
      6'b100101 : begin
        _zz_shift_q_6_6 = shift_q_map_37;
      end
      6'b100110 : begin
        _zz_shift_q_6_6 = shift_q_map_38;
      end
      default : begin
        _zz_shift_q_6_6 = shift_q_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_7_7)
      6'b000000 : begin
        _zz_shift_i_7_6 = shift_i_map_0;
      end
      6'b000001 : begin
        _zz_shift_i_7_6 = shift_i_map_1;
      end
      6'b000010 : begin
        _zz_shift_i_7_6 = shift_i_map_2;
      end
      6'b000011 : begin
        _zz_shift_i_7_6 = shift_i_map_3;
      end
      6'b000100 : begin
        _zz_shift_i_7_6 = shift_i_map_4;
      end
      6'b000101 : begin
        _zz_shift_i_7_6 = shift_i_map_5;
      end
      6'b000110 : begin
        _zz_shift_i_7_6 = shift_i_map_6;
      end
      6'b000111 : begin
        _zz_shift_i_7_6 = shift_i_map_7;
      end
      6'b001000 : begin
        _zz_shift_i_7_6 = shift_i_map_8;
      end
      6'b001001 : begin
        _zz_shift_i_7_6 = shift_i_map_9;
      end
      6'b001010 : begin
        _zz_shift_i_7_6 = shift_i_map_10;
      end
      6'b001011 : begin
        _zz_shift_i_7_6 = shift_i_map_11;
      end
      6'b001100 : begin
        _zz_shift_i_7_6 = shift_i_map_12;
      end
      6'b001101 : begin
        _zz_shift_i_7_6 = shift_i_map_13;
      end
      6'b001110 : begin
        _zz_shift_i_7_6 = shift_i_map_14;
      end
      6'b001111 : begin
        _zz_shift_i_7_6 = shift_i_map_15;
      end
      6'b010000 : begin
        _zz_shift_i_7_6 = shift_i_map_16;
      end
      6'b010001 : begin
        _zz_shift_i_7_6 = shift_i_map_17;
      end
      6'b010010 : begin
        _zz_shift_i_7_6 = shift_i_map_18;
      end
      6'b010011 : begin
        _zz_shift_i_7_6 = shift_i_map_19;
      end
      6'b010100 : begin
        _zz_shift_i_7_6 = shift_i_map_20;
      end
      6'b010101 : begin
        _zz_shift_i_7_6 = shift_i_map_21;
      end
      6'b010110 : begin
        _zz_shift_i_7_6 = shift_i_map_22;
      end
      6'b010111 : begin
        _zz_shift_i_7_6 = shift_i_map_23;
      end
      6'b011000 : begin
        _zz_shift_i_7_6 = shift_i_map_24;
      end
      6'b011001 : begin
        _zz_shift_i_7_6 = shift_i_map_25;
      end
      6'b011010 : begin
        _zz_shift_i_7_6 = shift_i_map_26;
      end
      6'b011011 : begin
        _zz_shift_i_7_6 = shift_i_map_27;
      end
      6'b011100 : begin
        _zz_shift_i_7_6 = shift_i_map_28;
      end
      6'b011101 : begin
        _zz_shift_i_7_6 = shift_i_map_29;
      end
      6'b011110 : begin
        _zz_shift_i_7_6 = shift_i_map_30;
      end
      6'b011111 : begin
        _zz_shift_i_7_6 = shift_i_map_31;
      end
      6'b100000 : begin
        _zz_shift_i_7_6 = shift_i_map_32;
      end
      6'b100001 : begin
        _zz_shift_i_7_6 = shift_i_map_33;
      end
      6'b100010 : begin
        _zz_shift_i_7_6 = shift_i_map_34;
      end
      6'b100011 : begin
        _zz_shift_i_7_6 = shift_i_map_35;
      end
      6'b100100 : begin
        _zz_shift_i_7_6 = shift_i_map_36;
      end
      6'b100101 : begin
        _zz_shift_i_7_6 = shift_i_map_37;
      end
      6'b100110 : begin
        _zz_shift_i_7_6 = shift_i_map_38;
      end
      default : begin
        _zz_shift_i_7_6 = shift_i_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_7_7)
      6'b000000 : begin
        _zz_shift_q_7_6 = shift_q_map_0;
      end
      6'b000001 : begin
        _zz_shift_q_7_6 = shift_q_map_1;
      end
      6'b000010 : begin
        _zz_shift_q_7_6 = shift_q_map_2;
      end
      6'b000011 : begin
        _zz_shift_q_7_6 = shift_q_map_3;
      end
      6'b000100 : begin
        _zz_shift_q_7_6 = shift_q_map_4;
      end
      6'b000101 : begin
        _zz_shift_q_7_6 = shift_q_map_5;
      end
      6'b000110 : begin
        _zz_shift_q_7_6 = shift_q_map_6;
      end
      6'b000111 : begin
        _zz_shift_q_7_6 = shift_q_map_7;
      end
      6'b001000 : begin
        _zz_shift_q_7_6 = shift_q_map_8;
      end
      6'b001001 : begin
        _zz_shift_q_7_6 = shift_q_map_9;
      end
      6'b001010 : begin
        _zz_shift_q_7_6 = shift_q_map_10;
      end
      6'b001011 : begin
        _zz_shift_q_7_6 = shift_q_map_11;
      end
      6'b001100 : begin
        _zz_shift_q_7_6 = shift_q_map_12;
      end
      6'b001101 : begin
        _zz_shift_q_7_6 = shift_q_map_13;
      end
      6'b001110 : begin
        _zz_shift_q_7_6 = shift_q_map_14;
      end
      6'b001111 : begin
        _zz_shift_q_7_6 = shift_q_map_15;
      end
      6'b010000 : begin
        _zz_shift_q_7_6 = shift_q_map_16;
      end
      6'b010001 : begin
        _zz_shift_q_7_6 = shift_q_map_17;
      end
      6'b010010 : begin
        _zz_shift_q_7_6 = shift_q_map_18;
      end
      6'b010011 : begin
        _zz_shift_q_7_6 = shift_q_map_19;
      end
      6'b010100 : begin
        _zz_shift_q_7_6 = shift_q_map_20;
      end
      6'b010101 : begin
        _zz_shift_q_7_6 = shift_q_map_21;
      end
      6'b010110 : begin
        _zz_shift_q_7_6 = shift_q_map_22;
      end
      6'b010111 : begin
        _zz_shift_q_7_6 = shift_q_map_23;
      end
      6'b011000 : begin
        _zz_shift_q_7_6 = shift_q_map_24;
      end
      6'b011001 : begin
        _zz_shift_q_7_6 = shift_q_map_25;
      end
      6'b011010 : begin
        _zz_shift_q_7_6 = shift_q_map_26;
      end
      6'b011011 : begin
        _zz_shift_q_7_6 = shift_q_map_27;
      end
      6'b011100 : begin
        _zz_shift_q_7_6 = shift_q_map_28;
      end
      6'b011101 : begin
        _zz_shift_q_7_6 = shift_q_map_29;
      end
      6'b011110 : begin
        _zz_shift_q_7_6 = shift_q_map_30;
      end
      6'b011111 : begin
        _zz_shift_q_7_6 = shift_q_map_31;
      end
      6'b100000 : begin
        _zz_shift_q_7_6 = shift_q_map_32;
      end
      6'b100001 : begin
        _zz_shift_q_7_6 = shift_q_map_33;
      end
      6'b100010 : begin
        _zz_shift_q_7_6 = shift_q_map_34;
      end
      6'b100011 : begin
        _zz_shift_q_7_6 = shift_q_map_35;
      end
      6'b100100 : begin
        _zz_shift_q_7_6 = shift_q_map_36;
      end
      6'b100101 : begin
        _zz_shift_q_7_6 = shift_q_map_37;
      end
      6'b100110 : begin
        _zz_shift_q_7_6 = shift_q_map_38;
      end
      default : begin
        _zz_shift_q_7_6 = shift_q_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_0_9)
      6'b000000 : begin
        _zz_shift_i_0_8 = shift_i_map_0;
      end
      6'b000001 : begin
        _zz_shift_i_0_8 = shift_i_map_1;
      end
      6'b000010 : begin
        _zz_shift_i_0_8 = shift_i_map_2;
      end
      6'b000011 : begin
        _zz_shift_i_0_8 = shift_i_map_3;
      end
      6'b000100 : begin
        _zz_shift_i_0_8 = shift_i_map_4;
      end
      6'b000101 : begin
        _zz_shift_i_0_8 = shift_i_map_5;
      end
      6'b000110 : begin
        _zz_shift_i_0_8 = shift_i_map_6;
      end
      6'b000111 : begin
        _zz_shift_i_0_8 = shift_i_map_7;
      end
      6'b001000 : begin
        _zz_shift_i_0_8 = shift_i_map_8;
      end
      6'b001001 : begin
        _zz_shift_i_0_8 = shift_i_map_9;
      end
      6'b001010 : begin
        _zz_shift_i_0_8 = shift_i_map_10;
      end
      6'b001011 : begin
        _zz_shift_i_0_8 = shift_i_map_11;
      end
      6'b001100 : begin
        _zz_shift_i_0_8 = shift_i_map_12;
      end
      6'b001101 : begin
        _zz_shift_i_0_8 = shift_i_map_13;
      end
      6'b001110 : begin
        _zz_shift_i_0_8 = shift_i_map_14;
      end
      6'b001111 : begin
        _zz_shift_i_0_8 = shift_i_map_15;
      end
      6'b010000 : begin
        _zz_shift_i_0_8 = shift_i_map_16;
      end
      6'b010001 : begin
        _zz_shift_i_0_8 = shift_i_map_17;
      end
      6'b010010 : begin
        _zz_shift_i_0_8 = shift_i_map_18;
      end
      6'b010011 : begin
        _zz_shift_i_0_8 = shift_i_map_19;
      end
      6'b010100 : begin
        _zz_shift_i_0_8 = shift_i_map_20;
      end
      6'b010101 : begin
        _zz_shift_i_0_8 = shift_i_map_21;
      end
      6'b010110 : begin
        _zz_shift_i_0_8 = shift_i_map_22;
      end
      6'b010111 : begin
        _zz_shift_i_0_8 = shift_i_map_23;
      end
      6'b011000 : begin
        _zz_shift_i_0_8 = shift_i_map_24;
      end
      6'b011001 : begin
        _zz_shift_i_0_8 = shift_i_map_25;
      end
      6'b011010 : begin
        _zz_shift_i_0_8 = shift_i_map_26;
      end
      6'b011011 : begin
        _zz_shift_i_0_8 = shift_i_map_27;
      end
      6'b011100 : begin
        _zz_shift_i_0_8 = shift_i_map_28;
      end
      6'b011101 : begin
        _zz_shift_i_0_8 = shift_i_map_29;
      end
      6'b011110 : begin
        _zz_shift_i_0_8 = shift_i_map_30;
      end
      6'b011111 : begin
        _zz_shift_i_0_8 = shift_i_map_31;
      end
      6'b100000 : begin
        _zz_shift_i_0_8 = shift_i_map_32;
      end
      6'b100001 : begin
        _zz_shift_i_0_8 = shift_i_map_33;
      end
      6'b100010 : begin
        _zz_shift_i_0_8 = shift_i_map_34;
      end
      6'b100011 : begin
        _zz_shift_i_0_8 = shift_i_map_35;
      end
      6'b100100 : begin
        _zz_shift_i_0_8 = shift_i_map_36;
      end
      6'b100101 : begin
        _zz_shift_i_0_8 = shift_i_map_37;
      end
      6'b100110 : begin
        _zz_shift_i_0_8 = shift_i_map_38;
      end
      default : begin
        _zz_shift_i_0_8 = shift_i_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_0_9)
      6'b000000 : begin
        _zz_shift_q_0_8 = shift_q_map_0;
      end
      6'b000001 : begin
        _zz_shift_q_0_8 = shift_q_map_1;
      end
      6'b000010 : begin
        _zz_shift_q_0_8 = shift_q_map_2;
      end
      6'b000011 : begin
        _zz_shift_q_0_8 = shift_q_map_3;
      end
      6'b000100 : begin
        _zz_shift_q_0_8 = shift_q_map_4;
      end
      6'b000101 : begin
        _zz_shift_q_0_8 = shift_q_map_5;
      end
      6'b000110 : begin
        _zz_shift_q_0_8 = shift_q_map_6;
      end
      6'b000111 : begin
        _zz_shift_q_0_8 = shift_q_map_7;
      end
      6'b001000 : begin
        _zz_shift_q_0_8 = shift_q_map_8;
      end
      6'b001001 : begin
        _zz_shift_q_0_8 = shift_q_map_9;
      end
      6'b001010 : begin
        _zz_shift_q_0_8 = shift_q_map_10;
      end
      6'b001011 : begin
        _zz_shift_q_0_8 = shift_q_map_11;
      end
      6'b001100 : begin
        _zz_shift_q_0_8 = shift_q_map_12;
      end
      6'b001101 : begin
        _zz_shift_q_0_8 = shift_q_map_13;
      end
      6'b001110 : begin
        _zz_shift_q_0_8 = shift_q_map_14;
      end
      6'b001111 : begin
        _zz_shift_q_0_8 = shift_q_map_15;
      end
      6'b010000 : begin
        _zz_shift_q_0_8 = shift_q_map_16;
      end
      6'b010001 : begin
        _zz_shift_q_0_8 = shift_q_map_17;
      end
      6'b010010 : begin
        _zz_shift_q_0_8 = shift_q_map_18;
      end
      6'b010011 : begin
        _zz_shift_q_0_8 = shift_q_map_19;
      end
      6'b010100 : begin
        _zz_shift_q_0_8 = shift_q_map_20;
      end
      6'b010101 : begin
        _zz_shift_q_0_8 = shift_q_map_21;
      end
      6'b010110 : begin
        _zz_shift_q_0_8 = shift_q_map_22;
      end
      6'b010111 : begin
        _zz_shift_q_0_8 = shift_q_map_23;
      end
      6'b011000 : begin
        _zz_shift_q_0_8 = shift_q_map_24;
      end
      6'b011001 : begin
        _zz_shift_q_0_8 = shift_q_map_25;
      end
      6'b011010 : begin
        _zz_shift_q_0_8 = shift_q_map_26;
      end
      6'b011011 : begin
        _zz_shift_q_0_8 = shift_q_map_27;
      end
      6'b011100 : begin
        _zz_shift_q_0_8 = shift_q_map_28;
      end
      6'b011101 : begin
        _zz_shift_q_0_8 = shift_q_map_29;
      end
      6'b011110 : begin
        _zz_shift_q_0_8 = shift_q_map_30;
      end
      6'b011111 : begin
        _zz_shift_q_0_8 = shift_q_map_31;
      end
      6'b100000 : begin
        _zz_shift_q_0_8 = shift_q_map_32;
      end
      6'b100001 : begin
        _zz_shift_q_0_8 = shift_q_map_33;
      end
      6'b100010 : begin
        _zz_shift_q_0_8 = shift_q_map_34;
      end
      6'b100011 : begin
        _zz_shift_q_0_8 = shift_q_map_35;
      end
      6'b100100 : begin
        _zz_shift_q_0_8 = shift_q_map_36;
      end
      6'b100101 : begin
        _zz_shift_q_0_8 = shift_q_map_37;
      end
      6'b100110 : begin
        _zz_shift_q_0_8 = shift_q_map_38;
      end
      default : begin
        _zz_shift_q_0_8 = shift_q_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_1_9)
      6'b000000 : begin
        _zz_shift_i_1_8 = shift_i_map_0;
      end
      6'b000001 : begin
        _zz_shift_i_1_8 = shift_i_map_1;
      end
      6'b000010 : begin
        _zz_shift_i_1_8 = shift_i_map_2;
      end
      6'b000011 : begin
        _zz_shift_i_1_8 = shift_i_map_3;
      end
      6'b000100 : begin
        _zz_shift_i_1_8 = shift_i_map_4;
      end
      6'b000101 : begin
        _zz_shift_i_1_8 = shift_i_map_5;
      end
      6'b000110 : begin
        _zz_shift_i_1_8 = shift_i_map_6;
      end
      6'b000111 : begin
        _zz_shift_i_1_8 = shift_i_map_7;
      end
      6'b001000 : begin
        _zz_shift_i_1_8 = shift_i_map_8;
      end
      6'b001001 : begin
        _zz_shift_i_1_8 = shift_i_map_9;
      end
      6'b001010 : begin
        _zz_shift_i_1_8 = shift_i_map_10;
      end
      6'b001011 : begin
        _zz_shift_i_1_8 = shift_i_map_11;
      end
      6'b001100 : begin
        _zz_shift_i_1_8 = shift_i_map_12;
      end
      6'b001101 : begin
        _zz_shift_i_1_8 = shift_i_map_13;
      end
      6'b001110 : begin
        _zz_shift_i_1_8 = shift_i_map_14;
      end
      6'b001111 : begin
        _zz_shift_i_1_8 = shift_i_map_15;
      end
      6'b010000 : begin
        _zz_shift_i_1_8 = shift_i_map_16;
      end
      6'b010001 : begin
        _zz_shift_i_1_8 = shift_i_map_17;
      end
      6'b010010 : begin
        _zz_shift_i_1_8 = shift_i_map_18;
      end
      6'b010011 : begin
        _zz_shift_i_1_8 = shift_i_map_19;
      end
      6'b010100 : begin
        _zz_shift_i_1_8 = shift_i_map_20;
      end
      6'b010101 : begin
        _zz_shift_i_1_8 = shift_i_map_21;
      end
      6'b010110 : begin
        _zz_shift_i_1_8 = shift_i_map_22;
      end
      6'b010111 : begin
        _zz_shift_i_1_8 = shift_i_map_23;
      end
      6'b011000 : begin
        _zz_shift_i_1_8 = shift_i_map_24;
      end
      6'b011001 : begin
        _zz_shift_i_1_8 = shift_i_map_25;
      end
      6'b011010 : begin
        _zz_shift_i_1_8 = shift_i_map_26;
      end
      6'b011011 : begin
        _zz_shift_i_1_8 = shift_i_map_27;
      end
      6'b011100 : begin
        _zz_shift_i_1_8 = shift_i_map_28;
      end
      6'b011101 : begin
        _zz_shift_i_1_8 = shift_i_map_29;
      end
      6'b011110 : begin
        _zz_shift_i_1_8 = shift_i_map_30;
      end
      6'b011111 : begin
        _zz_shift_i_1_8 = shift_i_map_31;
      end
      6'b100000 : begin
        _zz_shift_i_1_8 = shift_i_map_32;
      end
      6'b100001 : begin
        _zz_shift_i_1_8 = shift_i_map_33;
      end
      6'b100010 : begin
        _zz_shift_i_1_8 = shift_i_map_34;
      end
      6'b100011 : begin
        _zz_shift_i_1_8 = shift_i_map_35;
      end
      6'b100100 : begin
        _zz_shift_i_1_8 = shift_i_map_36;
      end
      6'b100101 : begin
        _zz_shift_i_1_8 = shift_i_map_37;
      end
      6'b100110 : begin
        _zz_shift_i_1_8 = shift_i_map_38;
      end
      default : begin
        _zz_shift_i_1_8 = shift_i_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_1_9)
      6'b000000 : begin
        _zz_shift_q_1_8 = shift_q_map_0;
      end
      6'b000001 : begin
        _zz_shift_q_1_8 = shift_q_map_1;
      end
      6'b000010 : begin
        _zz_shift_q_1_8 = shift_q_map_2;
      end
      6'b000011 : begin
        _zz_shift_q_1_8 = shift_q_map_3;
      end
      6'b000100 : begin
        _zz_shift_q_1_8 = shift_q_map_4;
      end
      6'b000101 : begin
        _zz_shift_q_1_8 = shift_q_map_5;
      end
      6'b000110 : begin
        _zz_shift_q_1_8 = shift_q_map_6;
      end
      6'b000111 : begin
        _zz_shift_q_1_8 = shift_q_map_7;
      end
      6'b001000 : begin
        _zz_shift_q_1_8 = shift_q_map_8;
      end
      6'b001001 : begin
        _zz_shift_q_1_8 = shift_q_map_9;
      end
      6'b001010 : begin
        _zz_shift_q_1_8 = shift_q_map_10;
      end
      6'b001011 : begin
        _zz_shift_q_1_8 = shift_q_map_11;
      end
      6'b001100 : begin
        _zz_shift_q_1_8 = shift_q_map_12;
      end
      6'b001101 : begin
        _zz_shift_q_1_8 = shift_q_map_13;
      end
      6'b001110 : begin
        _zz_shift_q_1_8 = shift_q_map_14;
      end
      6'b001111 : begin
        _zz_shift_q_1_8 = shift_q_map_15;
      end
      6'b010000 : begin
        _zz_shift_q_1_8 = shift_q_map_16;
      end
      6'b010001 : begin
        _zz_shift_q_1_8 = shift_q_map_17;
      end
      6'b010010 : begin
        _zz_shift_q_1_8 = shift_q_map_18;
      end
      6'b010011 : begin
        _zz_shift_q_1_8 = shift_q_map_19;
      end
      6'b010100 : begin
        _zz_shift_q_1_8 = shift_q_map_20;
      end
      6'b010101 : begin
        _zz_shift_q_1_8 = shift_q_map_21;
      end
      6'b010110 : begin
        _zz_shift_q_1_8 = shift_q_map_22;
      end
      6'b010111 : begin
        _zz_shift_q_1_8 = shift_q_map_23;
      end
      6'b011000 : begin
        _zz_shift_q_1_8 = shift_q_map_24;
      end
      6'b011001 : begin
        _zz_shift_q_1_8 = shift_q_map_25;
      end
      6'b011010 : begin
        _zz_shift_q_1_8 = shift_q_map_26;
      end
      6'b011011 : begin
        _zz_shift_q_1_8 = shift_q_map_27;
      end
      6'b011100 : begin
        _zz_shift_q_1_8 = shift_q_map_28;
      end
      6'b011101 : begin
        _zz_shift_q_1_8 = shift_q_map_29;
      end
      6'b011110 : begin
        _zz_shift_q_1_8 = shift_q_map_30;
      end
      6'b011111 : begin
        _zz_shift_q_1_8 = shift_q_map_31;
      end
      6'b100000 : begin
        _zz_shift_q_1_8 = shift_q_map_32;
      end
      6'b100001 : begin
        _zz_shift_q_1_8 = shift_q_map_33;
      end
      6'b100010 : begin
        _zz_shift_q_1_8 = shift_q_map_34;
      end
      6'b100011 : begin
        _zz_shift_q_1_8 = shift_q_map_35;
      end
      6'b100100 : begin
        _zz_shift_q_1_8 = shift_q_map_36;
      end
      6'b100101 : begin
        _zz_shift_q_1_8 = shift_q_map_37;
      end
      6'b100110 : begin
        _zz_shift_q_1_8 = shift_q_map_38;
      end
      default : begin
        _zz_shift_q_1_8 = shift_q_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_2_9)
      6'b000000 : begin
        _zz_shift_i_2_8 = shift_i_map_0;
      end
      6'b000001 : begin
        _zz_shift_i_2_8 = shift_i_map_1;
      end
      6'b000010 : begin
        _zz_shift_i_2_8 = shift_i_map_2;
      end
      6'b000011 : begin
        _zz_shift_i_2_8 = shift_i_map_3;
      end
      6'b000100 : begin
        _zz_shift_i_2_8 = shift_i_map_4;
      end
      6'b000101 : begin
        _zz_shift_i_2_8 = shift_i_map_5;
      end
      6'b000110 : begin
        _zz_shift_i_2_8 = shift_i_map_6;
      end
      6'b000111 : begin
        _zz_shift_i_2_8 = shift_i_map_7;
      end
      6'b001000 : begin
        _zz_shift_i_2_8 = shift_i_map_8;
      end
      6'b001001 : begin
        _zz_shift_i_2_8 = shift_i_map_9;
      end
      6'b001010 : begin
        _zz_shift_i_2_8 = shift_i_map_10;
      end
      6'b001011 : begin
        _zz_shift_i_2_8 = shift_i_map_11;
      end
      6'b001100 : begin
        _zz_shift_i_2_8 = shift_i_map_12;
      end
      6'b001101 : begin
        _zz_shift_i_2_8 = shift_i_map_13;
      end
      6'b001110 : begin
        _zz_shift_i_2_8 = shift_i_map_14;
      end
      6'b001111 : begin
        _zz_shift_i_2_8 = shift_i_map_15;
      end
      6'b010000 : begin
        _zz_shift_i_2_8 = shift_i_map_16;
      end
      6'b010001 : begin
        _zz_shift_i_2_8 = shift_i_map_17;
      end
      6'b010010 : begin
        _zz_shift_i_2_8 = shift_i_map_18;
      end
      6'b010011 : begin
        _zz_shift_i_2_8 = shift_i_map_19;
      end
      6'b010100 : begin
        _zz_shift_i_2_8 = shift_i_map_20;
      end
      6'b010101 : begin
        _zz_shift_i_2_8 = shift_i_map_21;
      end
      6'b010110 : begin
        _zz_shift_i_2_8 = shift_i_map_22;
      end
      6'b010111 : begin
        _zz_shift_i_2_8 = shift_i_map_23;
      end
      6'b011000 : begin
        _zz_shift_i_2_8 = shift_i_map_24;
      end
      6'b011001 : begin
        _zz_shift_i_2_8 = shift_i_map_25;
      end
      6'b011010 : begin
        _zz_shift_i_2_8 = shift_i_map_26;
      end
      6'b011011 : begin
        _zz_shift_i_2_8 = shift_i_map_27;
      end
      6'b011100 : begin
        _zz_shift_i_2_8 = shift_i_map_28;
      end
      6'b011101 : begin
        _zz_shift_i_2_8 = shift_i_map_29;
      end
      6'b011110 : begin
        _zz_shift_i_2_8 = shift_i_map_30;
      end
      6'b011111 : begin
        _zz_shift_i_2_8 = shift_i_map_31;
      end
      6'b100000 : begin
        _zz_shift_i_2_8 = shift_i_map_32;
      end
      6'b100001 : begin
        _zz_shift_i_2_8 = shift_i_map_33;
      end
      6'b100010 : begin
        _zz_shift_i_2_8 = shift_i_map_34;
      end
      6'b100011 : begin
        _zz_shift_i_2_8 = shift_i_map_35;
      end
      6'b100100 : begin
        _zz_shift_i_2_8 = shift_i_map_36;
      end
      6'b100101 : begin
        _zz_shift_i_2_8 = shift_i_map_37;
      end
      6'b100110 : begin
        _zz_shift_i_2_8 = shift_i_map_38;
      end
      default : begin
        _zz_shift_i_2_8 = shift_i_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_2_9)
      6'b000000 : begin
        _zz_shift_q_2_8 = shift_q_map_0;
      end
      6'b000001 : begin
        _zz_shift_q_2_8 = shift_q_map_1;
      end
      6'b000010 : begin
        _zz_shift_q_2_8 = shift_q_map_2;
      end
      6'b000011 : begin
        _zz_shift_q_2_8 = shift_q_map_3;
      end
      6'b000100 : begin
        _zz_shift_q_2_8 = shift_q_map_4;
      end
      6'b000101 : begin
        _zz_shift_q_2_8 = shift_q_map_5;
      end
      6'b000110 : begin
        _zz_shift_q_2_8 = shift_q_map_6;
      end
      6'b000111 : begin
        _zz_shift_q_2_8 = shift_q_map_7;
      end
      6'b001000 : begin
        _zz_shift_q_2_8 = shift_q_map_8;
      end
      6'b001001 : begin
        _zz_shift_q_2_8 = shift_q_map_9;
      end
      6'b001010 : begin
        _zz_shift_q_2_8 = shift_q_map_10;
      end
      6'b001011 : begin
        _zz_shift_q_2_8 = shift_q_map_11;
      end
      6'b001100 : begin
        _zz_shift_q_2_8 = shift_q_map_12;
      end
      6'b001101 : begin
        _zz_shift_q_2_8 = shift_q_map_13;
      end
      6'b001110 : begin
        _zz_shift_q_2_8 = shift_q_map_14;
      end
      6'b001111 : begin
        _zz_shift_q_2_8 = shift_q_map_15;
      end
      6'b010000 : begin
        _zz_shift_q_2_8 = shift_q_map_16;
      end
      6'b010001 : begin
        _zz_shift_q_2_8 = shift_q_map_17;
      end
      6'b010010 : begin
        _zz_shift_q_2_8 = shift_q_map_18;
      end
      6'b010011 : begin
        _zz_shift_q_2_8 = shift_q_map_19;
      end
      6'b010100 : begin
        _zz_shift_q_2_8 = shift_q_map_20;
      end
      6'b010101 : begin
        _zz_shift_q_2_8 = shift_q_map_21;
      end
      6'b010110 : begin
        _zz_shift_q_2_8 = shift_q_map_22;
      end
      6'b010111 : begin
        _zz_shift_q_2_8 = shift_q_map_23;
      end
      6'b011000 : begin
        _zz_shift_q_2_8 = shift_q_map_24;
      end
      6'b011001 : begin
        _zz_shift_q_2_8 = shift_q_map_25;
      end
      6'b011010 : begin
        _zz_shift_q_2_8 = shift_q_map_26;
      end
      6'b011011 : begin
        _zz_shift_q_2_8 = shift_q_map_27;
      end
      6'b011100 : begin
        _zz_shift_q_2_8 = shift_q_map_28;
      end
      6'b011101 : begin
        _zz_shift_q_2_8 = shift_q_map_29;
      end
      6'b011110 : begin
        _zz_shift_q_2_8 = shift_q_map_30;
      end
      6'b011111 : begin
        _zz_shift_q_2_8 = shift_q_map_31;
      end
      6'b100000 : begin
        _zz_shift_q_2_8 = shift_q_map_32;
      end
      6'b100001 : begin
        _zz_shift_q_2_8 = shift_q_map_33;
      end
      6'b100010 : begin
        _zz_shift_q_2_8 = shift_q_map_34;
      end
      6'b100011 : begin
        _zz_shift_q_2_8 = shift_q_map_35;
      end
      6'b100100 : begin
        _zz_shift_q_2_8 = shift_q_map_36;
      end
      6'b100101 : begin
        _zz_shift_q_2_8 = shift_q_map_37;
      end
      6'b100110 : begin
        _zz_shift_q_2_8 = shift_q_map_38;
      end
      default : begin
        _zz_shift_q_2_8 = shift_q_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_3_9)
      6'b000000 : begin
        _zz_shift_i_3_8 = shift_i_map_0;
      end
      6'b000001 : begin
        _zz_shift_i_3_8 = shift_i_map_1;
      end
      6'b000010 : begin
        _zz_shift_i_3_8 = shift_i_map_2;
      end
      6'b000011 : begin
        _zz_shift_i_3_8 = shift_i_map_3;
      end
      6'b000100 : begin
        _zz_shift_i_3_8 = shift_i_map_4;
      end
      6'b000101 : begin
        _zz_shift_i_3_8 = shift_i_map_5;
      end
      6'b000110 : begin
        _zz_shift_i_3_8 = shift_i_map_6;
      end
      6'b000111 : begin
        _zz_shift_i_3_8 = shift_i_map_7;
      end
      6'b001000 : begin
        _zz_shift_i_3_8 = shift_i_map_8;
      end
      6'b001001 : begin
        _zz_shift_i_3_8 = shift_i_map_9;
      end
      6'b001010 : begin
        _zz_shift_i_3_8 = shift_i_map_10;
      end
      6'b001011 : begin
        _zz_shift_i_3_8 = shift_i_map_11;
      end
      6'b001100 : begin
        _zz_shift_i_3_8 = shift_i_map_12;
      end
      6'b001101 : begin
        _zz_shift_i_3_8 = shift_i_map_13;
      end
      6'b001110 : begin
        _zz_shift_i_3_8 = shift_i_map_14;
      end
      6'b001111 : begin
        _zz_shift_i_3_8 = shift_i_map_15;
      end
      6'b010000 : begin
        _zz_shift_i_3_8 = shift_i_map_16;
      end
      6'b010001 : begin
        _zz_shift_i_3_8 = shift_i_map_17;
      end
      6'b010010 : begin
        _zz_shift_i_3_8 = shift_i_map_18;
      end
      6'b010011 : begin
        _zz_shift_i_3_8 = shift_i_map_19;
      end
      6'b010100 : begin
        _zz_shift_i_3_8 = shift_i_map_20;
      end
      6'b010101 : begin
        _zz_shift_i_3_8 = shift_i_map_21;
      end
      6'b010110 : begin
        _zz_shift_i_3_8 = shift_i_map_22;
      end
      6'b010111 : begin
        _zz_shift_i_3_8 = shift_i_map_23;
      end
      6'b011000 : begin
        _zz_shift_i_3_8 = shift_i_map_24;
      end
      6'b011001 : begin
        _zz_shift_i_3_8 = shift_i_map_25;
      end
      6'b011010 : begin
        _zz_shift_i_3_8 = shift_i_map_26;
      end
      6'b011011 : begin
        _zz_shift_i_3_8 = shift_i_map_27;
      end
      6'b011100 : begin
        _zz_shift_i_3_8 = shift_i_map_28;
      end
      6'b011101 : begin
        _zz_shift_i_3_8 = shift_i_map_29;
      end
      6'b011110 : begin
        _zz_shift_i_3_8 = shift_i_map_30;
      end
      6'b011111 : begin
        _zz_shift_i_3_8 = shift_i_map_31;
      end
      6'b100000 : begin
        _zz_shift_i_3_8 = shift_i_map_32;
      end
      6'b100001 : begin
        _zz_shift_i_3_8 = shift_i_map_33;
      end
      6'b100010 : begin
        _zz_shift_i_3_8 = shift_i_map_34;
      end
      6'b100011 : begin
        _zz_shift_i_3_8 = shift_i_map_35;
      end
      6'b100100 : begin
        _zz_shift_i_3_8 = shift_i_map_36;
      end
      6'b100101 : begin
        _zz_shift_i_3_8 = shift_i_map_37;
      end
      6'b100110 : begin
        _zz_shift_i_3_8 = shift_i_map_38;
      end
      default : begin
        _zz_shift_i_3_8 = shift_i_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_3_9)
      6'b000000 : begin
        _zz_shift_q_3_8 = shift_q_map_0;
      end
      6'b000001 : begin
        _zz_shift_q_3_8 = shift_q_map_1;
      end
      6'b000010 : begin
        _zz_shift_q_3_8 = shift_q_map_2;
      end
      6'b000011 : begin
        _zz_shift_q_3_8 = shift_q_map_3;
      end
      6'b000100 : begin
        _zz_shift_q_3_8 = shift_q_map_4;
      end
      6'b000101 : begin
        _zz_shift_q_3_8 = shift_q_map_5;
      end
      6'b000110 : begin
        _zz_shift_q_3_8 = shift_q_map_6;
      end
      6'b000111 : begin
        _zz_shift_q_3_8 = shift_q_map_7;
      end
      6'b001000 : begin
        _zz_shift_q_3_8 = shift_q_map_8;
      end
      6'b001001 : begin
        _zz_shift_q_3_8 = shift_q_map_9;
      end
      6'b001010 : begin
        _zz_shift_q_3_8 = shift_q_map_10;
      end
      6'b001011 : begin
        _zz_shift_q_3_8 = shift_q_map_11;
      end
      6'b001100 : begin
        _zz_shift_q_3_8 = shift_q_map_12;
      end
      6'b001101 : begin
        _zz_shift_q_3_8 = shift_q_map_13;
      end
      6'b001110 : begin
        _zz_shift_q_3_8 = shift_q_map_14;
      end
      6'b001111 : begin
        _zz_shift_q_3_8 = shift_q_map_15;
      end
      6'b010000 : begin
        _zz_shift_q_3_8 = shift_q_map_16;
      end
      6'b010001 : begin
        _zz_shift_q_3_8 = shift_q_map_17;
      end
      6'b010010 : begin
        _zz_shift_q_3_8 = shift_q_map_18;
      end
      6'b010011 : begin
        _zz_shift_q_3_8 = shift_q_map_19;
      end
      6'b010100 : begin
        _zz_shift_q_3_8 = shift_q_map_20;
      end
      6'b010101 : begin
        _zz_shift_q_3_8 = shift_q_map_21;
      end
      6'b010110 : begin
        _zz_shift_q_3_8 = shift_q_map_22;
      end
      6'b010111 : begin
        _zz_shift_q_3_8 = shift_q_map_23;
      end
      6'b011000 : begin
        _zz_shift_q_3_8 = shift_q_map_24;
      end
      6'b011001 : begin
        _zz_shift_q_3_8 = shift_q_map_25;
      end
      6'b011010 : begin
        _zz_shift_q_3_8 = shift_q_map_26;
      end
      6'b011011 : begin
        _zz_shift_q_3_8 = shift_q_map_27;
      end
      6'b011100 : begin
        _zz_shift_q_3_8 = shift_q_map_28;
      end
      6'b011101 : begin
        _zz_shift_q_3_8 = shift_q_map_29;
      end
      6'b011110 : begin
        _zz_shift_q_3_8 = shift_q_map_30;
      end
      6'b011111 : begin
        _zz_shift_q_3_8 = shift_q_map_31;
      end
      6'b100000 : begin
        _zz_shift_q_3_8 = shift_q_map_32;
      end
      6'b100001 : begin
        _zz_shift_q_3_8 = shift_q_map_33;
      end
      6'b100010 : begin
        _zz_shift_q_3_8 = shift_q_map_34;
      end
      6'b100011 : begin
        _zz_shift_q_3_8 = shift_q_map_35;
      end
      6'b100100 : begin
        _zz_shift_q_3_8 = shift_q_map_36;
      end
      6'b100101 : begin
        _zz_shift_q_3_8 = shift_q_map_37;
      end
      6'b100110 : begin
        _zz_shift_q_3_8 = shift_q_map_38;
      end
      default : begin
        _zz_shift_q_3_8 = shift_q_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_4_9)
      6'b000000 : begin
        _zz_shift_i_4_8 = shift_i_map_0;
      end
      6'b000001 : begin
        _zz_shift_i_4_8 = shift_i_map_1;
      end
      6'b000010 : begin
        _zz_shift_i_4_8 = shift_i_map_2;
      end
      6'b000011 : begin
        _zz_shift_i_4_8 = shift_i_map_3;
      end
      6'b000100 : begin
        _zz_shift_i_4_8 = shift_i_map_4;
      end
      6'b000101 : begin
        _zz_shift_i_4_8 = shift_i_map_5;
      end
      6'b000110 : begin
        _zz_shift_i_4_8 = shift_i_map_6;
      end
      6'b000111 : begin
        _zz_shift_i_4_8 = shift_i_map_7;
      end
      6'b001000 : begin
        _zz_shift_i_4_8 = shift_i_map_8;
      end
      6'b001001 : begin
        _zz_shift_i_4_8 = shift_i_map_9;
      end
      6'b001010 : begin
        _zz_shift_i_4_8 = shift_i_map_10;
      end
      6'b001011 : begin
        _zz_shift_i_4_8 = shift_i_map_11;
      end
      6'b001100 : begin
        _zz_shift_i_4_8 = shift_i_map_12;
      end
      6'b001101 : begin
        _zz_shift_i_4_8 = shift_i_map_13;
      end
      6'b001110 : begin
        _zz_shift_i_4_8 = shift_i_map_14;
      end
      6'b001111 : begin
        _zz_shift_i_4_8 = shift_i_map_15;
      end
      6'b010000 : begin
        _zz_shift_i_4_8 = shift_i_map_16;
      end
      6'b010001 : begin
        _zz_shift_i_4_8 = shift_i_map_17;
      end
      6'b010010 : begin
        _zz_shift_i_4_8 = shift_i_map_18;
      end
      6'b010011 : begin
        _zz_shift_i_4_8 = shift_i_map_19;
      end
      6'b010100 : begin
        _zz_shift_i_4_8 = shift_i_map_20;
      end
      6'b010101 : begin
        _zz_shift_i_4_8 = shift_i_map_21;
      end
      6'b010110 : begin
        _zz_shift_i_4_8 = shift_i_map_22;
      end
      6'b010111 : begin
        _zz_shift_i_4_8 = shift_i_map_23;
      end
      6'b011000 : begin
        _zz_shift_i_4_8 = shift_i_map_24;
      end
      6'b011001 : begin
        _zz_shift_i_4_8 = shift_i_map_25;
      end
      6'b011010 : begin
        _zz_shift_i_4_8 = shift_i_map_26;
      end
      6'b011011 : begin
        _zz_shift_i_4_8 = shift_i_map_27;
      end
      6'b011100 : begin
        _zz_shift_i_4_8 = shift_i_map_28;
      end
      6'b011101 : begin
        _zz_shift_i_4_8 = shift_i_map_29;
      end
      6'b011110 : begin
        _zz_shift_i_4_8 = shift_i_map_30;
      end
      6'b011111 : begin
        _zz_shift_i_4_8 = shift_i_map_31;
      end
      6'b100000 : begin
        _zz_shift_i_4_8 = shift_i_map_32;
      end
      6'b100001 : begin
        _zz_shift_i_4_8 = shift_i_map_33;
      end
      6'b100010 : begin
        _zz_shift_i_4_8 = shift_i_map_34;
      end
      6'b100011 : begin
        _zz_shift_i_4_8 = shift_i_map_35;
      end
      6'b100100 : begin
        _zz_shift_i_4_8 = shift_i_map_36;
      end
      6'b100101 : begin
        _zz_shift_i_4_8 = shift_i_map_37;
      end
      6'b100110 : begin
        _zz_shift_i_4_8 = shift_i_map_38;
      end
      default : begin
        _zz_shift_i_4_8 = shift_i_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_4_9)
      6'b000000 : begin
        _zz_shift_q_4_8 = shift_q_map_0;
      end
      6'b000001 : begin
        _zz_shift_q_4_8 = shift_q_map_1;
      end
      6'b000010 : begin
        _zz_shift_q_4_8 = shift_q_map_2;
      end
      6'b000011 : begin
        _zz_shift_q_4_8 = shift_q_map_3;
      end
      6'b000100 : begin
        _zz_shift_q_4_8 = shift_q_map_4;
      end
      6'b000101 : begin
        _zz_shift_q_4_8 = shift_q_map_5;
      end
      6'b000110 : begin
        _zz_shift_q_4_8 = shift_q_map_6;
      end
      6'b000111 : begin
        _zz_shift_q_4_8 = shift_q_map_7;
      end
      6'b001000 : begin
        _zz_shift_q_4_8 = shift_q_map_8;
      end
      6'b001001 : begin
        _zz_shift_q_4_8 = shift_q_map_9;
      end
      6'b001010 : begin
        _zz_shift_q_4_8 = shift_q_map_10;
      end
      6'b001011 : begin
        _zz_shift_q_4_8 = shift_q_map_11;
      end
      6'b001100 : begin
        _zz_shift_q_4_8 = shift_q_map_12;
      end
      6'b001101 : begin
        _zz_shift_q_4_8 = shift_q_map_13;
      end
      6'b001110 : begin
        _zz_shift_q_4_8 = shift_q_map_14;
      end
      6'b001111 : begin
        _zz_shift_q_4_8 = shift_q_map_15;
      end
      6'b010000 : begin
        _zz_shift_q_4_8 = shift_q_map_16;
      end
      6'b010001 : begin
        _zz_shift_q_4_8 = shift_q_map_17;
      end
      6'b010010 : begin
        _zz_shift_q_4_8 = shift_q_map_18;
      end
      6'b010011 : begin
        _zz_shift_q_4_8 = shift_q_map_19;
      end
      6'b010100 : begin
        _zz_shift_q_4_8 = shift_q_map_20;
      end
      6'b010101 : begin
        _zz_shift_q_4_8 = shift_q_map_21;
      end
      6'b010110 : begin
        _zz_shift_q_4_8 = shift_q_map_22;
      end
      6'b010111 : begin
        _zz_shift_q_4_8 = shift_q_map_23;
      end
      6'b011000 : begin
        _zz_shift_q_4_8 = shift_q_map_24;
      end
      6'b011001 : begin
        _zz_shift_q_4_8 = shift_q_map_25;
      end
      6'b011010 : begin
        _zz_shift_q_4_8 = shift_q_map_26;
      end
      6'b011011 : begin
        _zz_shift_q_4_8 = shift_q_map_27;
      end
      6'b011100 : begin
        _zz_shift_q_4_8 = shift_q_map_28;
      end
      6'b011101 : begin
        _zz_shift_q_4_8 = shift_q_map_29;
      end
      6'b011110 : begin
        _zz_shift_q_4_8 = shift_q_map_30;
      end
      6'b011111 : begin
        _zz_shift_q_4_8 = shift_q_map_31;
      end
      6'b100000 : begin
        _zz_shift_q_4_8 = shift_q_map_32;
      end
      6'b100001 : begin
        _zz_shift_q_4_8 = shift_q_map_33;
      end
      6'b100010 : begin
        _zz_shift_q_4_8 = shift_q_map_34;
      end
      6'b100011 : begin
        _zz_shift_q_4_8 = shift_q_map_35;
      end
      6'b100100 : begin
        _zz_shift_q_4_8 = shift_q_map_36;
      end
      6'b100101 : begin
        _zz_shift_q_4_8 = shift_q_map_37;
      end
      6'b100110 : begin
        _zz_shift_q_4_8 = shift_q_map_38;
      end
      default : begin
        _zz_shift_q_4_8 = shift_q_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_5_9)
      6'b000000 : begin
        _zz_shift_i_5_8 = shift_i_map_0;
      end
      6'b000001 : begin
        _zz_shift_i_5_8 = shift_i_map_1;
      end
      6'b000010 : begin
        _zz_shift_i_5_8 = shift_i_map_2;
      end
      6'b000011 : begin
        _zz_shift_i_5_8 = shift_i_map_3;
      end
      6'b000100 : begin
        _zz_shift_i_5_8 = shift_i_map_4;
      end
      6'b000101 : begin
        _zz_shift_i_5_8 = shift_i_map_5;
      end
      6'b000110 : begin
        _zz_shift_i_5_8 = shift_i_map_6;
      end
      6'b000111 : begin
        _zz_shift_i_5_8 = shift_i_map_7;
      end
      6'b001000 : begin
        _zz_shift_i_5_8 = shift_i_map_8;
      end
      6'b001001 : begin
        _zz_shift_i_5_8 = shift_i_map_9;
      end
      6'b001010 : begin
        _zz_shift_i_5_8 = shift_i_map_10;
      end
      6'b001011 : begin
        _zz_shift_i_5_8 = shift_i_map_11;
      end
      6'b001100 : begin
        _zz_shift_i_5_8 = shift_i_map_12;
      end
      6'b001101 : begin
        _zz_shift_i_5_8 = shift_i_map_13;
      end
      6'b001110 : begin
        _zz_shift_i_5_8 = shift_i_map_14;
      end
      6'b001111 : begin
        _zz_shift_i_5_8 = shift_i_map_15;
      end
      6'b010000 : begin
        _zz_shift_i_5_8 = shift_i_map_16;
      end
      6'b010001 : begin
        _zz_shift_i_5_8 = shift_i_map_17;
      end
      6'b010010 : begin
        _zz_shift_i_5_8 = shift_i_map_18;
      end
      6'b010011 : begin
        _zz_shift_i_5_8 = shift_i_map_19;
      end
      6'b010100 : begin
        _zz_shift_i_5_8 = shift_i_map_20;
      end
      6'b010101 : begin
        _zz_shift_i_5_8 = shift_i_map_21;
      end
      6'b010110 : begin
        _zz_shift_i_5_8 = shift_i_map_22;
      end
      6'b010111 : begin
        _zz_shift_i_5_8 = shift_i_map_23;
      end
      6'b011000 : begin
        _zz_shift_i_5_8 = shift_i_map_24;
      end
      6'b011001 : begin
        _zz_shift_i_5_8 = shift_i_map_25;
      end
      6'b011010 : begin
        _zz_shift_i_5_8 = shift_i_map_26;
      end
      6'b011011 : begin
        _zz_shift_i_5_8 = shift_i_map_27;
      end
      6'b011100 : begin
        _zz_shift_i_5_8 = shift_i_map_28;
      end
      6'b011101 : begin
        _zz_shift_i_5_8 = shift_i_map_29;
      end
      6'b011110 : begin
        _zz_shift_i_5_8 = shift_i_map_30;
      end
      6'b011111 : begin
        _zz_shift_i_5_8 = shift_i_map_31;
      end
      6'b100000 : begin
        _zz_shift_i_5_8 = shift_i_map_32;
      end
      6'b100001 : begin
        _zz_shift_i_5_8 = shift_i_map_33;
      end
      6'b100010 : begin
        _zz_shift_i_5_8 = shift_i_map_34;
      end
      6'b100011 : begin
        _zz_shift_i_5_8 = shift_i_map_35;
      end
      6'b100100 : begin
        _zz_shift_i_5_8 = shift_i_map_36;
      end
      6'b100101 : begin
        _zz_shift_i_5_8 = shift_i_map_37;
      end
      6'b100110 : begin
        _zz_shift_i_5_8 = shift_i_map_38;
      end
      default : begin
        _zz_shift_i_5_8 = shift_i_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_5_9)
      6'b000000 : begin
        _zz_shift_q_5_8 = shift_q_map_0;
      end
      6'b000001 : begin
        _zz_shift_q_5_8 = shift_q_map_1;
      end
      6'b000010 : begin
        _zz_shift_q_5_8 = shift_q_map_2;
      end
      6'b000011 : begin
        _zz_shift_q_5_8 = shift_q_map_3;
      end
      6'b000100 : begin
        _zz_shift_q_5_8 = shift_q_map_4;
      end
      6'b000101 : begin
        _zz_shift_q_5_8 = shift_q_map_5;
      end
      6'b000110 : begin
        _zz_shift_q_5_8 = shift_q_map_6;
      end
      6'b000111 : begin
        _zz_shift_q_5_8 = shift_q_map_7;
      end
      6'b001000 : begin
        _zz_shift_q_5_8 = shift_q_map_8;
      end
      6'b001001 : begin
        _zz_shift_q_5_8 = shift_q_map_9;
      end
      6'b001010 : begin
        _zz_shift_q_5_8 = shift_q_map_10;
      end
      6'b001011 : begin
        _zz_shift_q_5_8 = shift_q_map_11;
      end
      6'b001100 : begin
        _zz_shift_q_5_8 = shift_q_map_12;
      end
      6'b001101 : begin
        _zz_shift_q_5_8 = shift_q_map_13;
      end
      6'b001110 : begin
        _zz_shift_q_5_8 = shift_q_map_14;
      end
      6'b001111 : begin
        _zz_shift_q_5_8 = shift_q_map_15;
      end
      6'b010000 : begin
        _zz_shift_q_5_8 = shift_q_map_16;
      end
      6'b010001 : begin
        _zz_shift_q_5_8 = shift_q_map_17;
      end
      6'b010010 : begin
        _zz_shift_q_5_8 = shift_q_map_18;
      end
      6'b010011 : begin
        _zz_shift_q_5_8 = shift_q_map_19;
      end
      6'b010100 : begin
        _zz_shift_q_5_8 = shift_q_map_20;
      end
      6'b010101 : begin
        _zz_shift_q_5_8 = shift_q_map_21;
      end
      6'b010110 : begin
        _zz_shift_q_5_8 = shift_q_map_22;
      end
      6'b010111 : begin
        _zz_shift_q_5_8 = shift_q_map_23;
      end
      6'b011000 : begin
        _zz_shift_q_5_8 = shift_q_map_24;
      end
      6'b011001 : begin
        _zz_shift_q_5_8 = shift_q_map_25;
      end
      6'b011010 : begin
        _zz_shift_q_5_8 = shift_q_map_26;
      end
      6'b011011 : begin
        _zz_shift_q_5_8 = shift_q_map_27;
      end
      6'b011100 : begin
        _zz_shift_q_5_8 = shift_q_map_28;
      end
      6'b011101 : begin
        _zz_shift_q_5_8 = shift_q_map_29;
      end
      6'b011110 : begin
        _zz_shift_q_5_8 = shift_q_map_30;
      end
      6'b011111 : begin
        _zz_shift_q_5_8 = shift_q_map_31;
      end
      6'b100000 : begin
        _zz_shift_q_5_8 = shift_q_map_32;
      end
      6'b100001 : begin
        _zz_shift_q_5_8 = shift_q_map_33;
      end
      6'b100010 : begin
        _zz_shift_q_5_8 = shift_q_map_34;
      end
      6'b100011 : begin
        _zz_shift_q_5_8 = shift_q_map_35;
      end
      6'b100100 : begin
        _zz_shift_q_5_8 = shift_q_map_36;
      end
      6'b100101 : begin
        _zz_shift_q_5_8 = shift_q_map_37;
      end
      6'b100110 : begin
        _zz_shift_q_5_8 = shift_q_map_38;
      end
      default : begin
        _zz_shift_q_5_8 = shift_q_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_6_9)
      6'b000000 : begin
        _zz_shift_i_6_8 = shift_i_map_0;
      end
      6'b000001 : begin
        _zz_shift_i_6_8 = shift_i_map_1;
      end
      6'b000010 : begin
        _zz_shift_i_6_8 = shift_i_map_2;
      end
      6'b000011 : begin
        _zz_shift_i_6_8 = shift_i_map_3;
      end
      6'b000100 : begin
        _zz_shift_i_6_8 = shift_i_map_4;
      end
      6'b000101 : begin
        _zz_shift_i_6_8 = shift_i_map_5;
      end
      6'b000110 : begin
        _zz_shift_i_6_8 = shift_i_map_6;
      end
      6'b000111 : begin
        _zz_shift_i_6_8 = shift_i_map_7;
      end
      6'b001000 : begin
        _zz_shift_i_6_8 = shift_i_map_8;
      end
      6'b001001 : begin
        _zz_shift_i_6_8 = shift_i_map_9;
      end
      6'b001010 : begin
        _zz_shift_i_6_8 = shift_i_map_10;
      end
      6'b001011 : begin
        _zz_shift_i_6_8 = shift_i_map_11;
      end
      6'b001100 : begin
        _zz_shift_i_6_8 = shift_i_map_12;
      end
      6'b001101 : begin
        _zz_shift_i_6_8 = shift_i_map_13;
      end
      6'b001110 : begin
        _zz_shift_i_6_8 = shift_i_map_14;
      end
      6'b001111 : begin
        _zz_shift_i_6_8 = shift_i_map_15;
      end
      6'b010000 : begin
        _zz_shift_i_6_8 = shift_i_map_16;
      end
      6'b010001 : begin
        _zz_shift_i_6_8 = shift_i_map_17;
      end
      6'b010010 : begin
        _zz_shift_i_6_8 = shift_i_map_18;
      end
      6'b010011 : begin
        _zz_shift_i_6_8 = shift_i_map_19;
      end
      6'b010100 : begin
        _zz_shift_i_6_8 = shift_i_map_20;
      end
      6'b010101 : begin
        _zz_shift_i_6_8 = shift_i_map_21;
      end
      6'b010110 : begin
        _zz_shift_i_6_8 = shift_i_map_22;
      end
      6'b010111 : begin
        _zz_shift_i_6_8 = shift_i_map_23;
      end
      6'b011000 : begin
        _zz_shift_i_6_8 = shift_i_map_24;
      end
      6'b011001 : begin
        _zz_shift_i_6_8 = shift_i_map_25;
      end
      6'b011010 : begin
        _zz_shift_i_6_8 = shift_i_map_26;
      end
      6'b011011 : begin
        _zz_shift_i_6_8 = shift_i_map_27;
      end
      6'b011100 : begin
        _zz_shift_i_6_8 = shift_i_map_28;
      end
      6'b011101 : begin
        _zz_shift_i_6_8 = shift_i_map_29;
      end
      6'b011110 : begin
        _zz_shift_i_6_8 = shift_i_map_30;
      end
      6'b011111 : begin
        _zz_shift_i_6_8 = shift_i_map_31;
      end
      6'b100000 : begin
        _zz_shift_i_6_8 = shift_i_map_32;
      end
      6'b100001 : begin
        _zz_shift_i_6_8 = shift_i_map_33;
      end
      6'b100010 : begin
        _zz_shift_i_6_8 = shift_i_map_34;
      end
      6'b100011 : begin
        _zz_shift_i_6_8 = shift_i_map_35;
      end
      6'b100100 : begin
        _zz_shift_i_6_8 = shift_i_map_36;
      end
      6'b100101 : begin
        _zz_shift_i_6_8 = shift_i_map_37;
      end
      6'b100110 : begin
        _zz_shift_i_6_8 = shift_i_map_38;
      end
      default : begin
        _zz_shift_i_6_8 = shift_i_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_6_9)
      6'b000000 : begin
        _zz_shift_q_6_8 = shift_q_map_0;
      end
      6'b000001 : begin
        _zz_shift_q_6_8 = shift_q_map_1;
      end
      6'b000010 : begin
        _zz_shift_q_6_8 = shift_q_map_2;
      end
      6'b000011 : begin
        _zz_shift_q_6_8 = shift_q_map_3;
      end
      6'b000100 : begin
        _zz_shift_q_6_8 = shift_q_map_4;
      end
      6'b000101 : begin
        _zz_shift_q_6_8 = shift_q_map_5;
      end
      6'b000110 : begin
        _zz_shift_q_6_8 = shift_q_map_6;
      end
      6'b000111 : begin
        _zz_shift_q_6_8 = shift_q_map_7;
      end
      6'b001000 : begin
        _zz_shift_q_6_8 = shift_q_map_8;
      end
      6'b001001 : begin
        _zz_shift_q_6_8 = shift_q_map_9;
      end
      6'b001010 : begin
        _zz_shift_q_6_8 = shift_q_map_10;
      end
      6'b001011 : begin
        _zz_shift_q_6_8 = shift_q_map_11;
      end
      6'b001100 : begin
        _zz_shift_q_6_8 = shift_q_map_12;
      end
      6'b001101 : begin
        _zz_shift_q_6_8 = shift_q_map_13;
      end
      6'b001110 : begin
        _zz_shift_q_6_8 = shift_q_map_14;
      end
      6'b001111 : begin
        _zz_shift_q_6_8 = shift_q_map_15;
      end
      6'b010000 : begin
        _zz_shift_q_6_8 = shift_q_map_16;
      end
      6'b010001 : begin
        _zz_shift_q_6_8 = shift_q_map_17;
      end
      6'b010010 : begin
        _zz_shift_q_6_8 = shift_q_map_18;
      end
      6'b010011 : begin
        _zz_shift_q_6_8 = shift_q_map_19;
      end
      6'b010100 : begin
        _zz_shift_q_6_8 = shift_q_map_20;
      end
      6'b010101 : begin
        _zz_shift_q_6_8 = shift_q_map_21;
      end
      6'b010110 : begin
        _zz_shift_q_6_8 = shift_q_map_22;
      end
      6'b010111 : begin
        _zz_shift_q_6_8 = shift_q_map_23;
      end
      6'b011000 : begin
        _zz_shift_q_6_8 = shift_q_map_24;
      end
      6'b011001 : begin
        _zz_shift_q_6_8 = shift_q_map_25;
      end
      6'b011010 : begin
        _zz_shift_q_6_8 = shift_q_map_26;
      end
      6'b011011 : begin
        _zz_shift_q_6_8 = shift_q_map_27;
      end
      6'b011100 : begin
        _zz_shift_q_6_8 = shift_q_map_28;
      end
      6'b011101 : begin
        _zz_shift_q_6_8 = shift_q_map_29;
      end
      6'b011110 : begin
        _zz_shift_q_6_8 = shift_q_map_30;
      end
      6'b011111 : begin
        _zz_shift_q_6_8 = shift_q_map_31;
      end
      6'b100000 : begin
        _zz_shift_q_6_8 = shift_q_map_32;
      end
      6'b100001 : begin
        _zz_shift_q_6_8 = shift_q_map_33;
      end
      6'b100010 : begin
        _zz_shift_q_6_8 = shift_q_map_34;
      end
      6'b100011 : begin
        _zz_shift_q_6_8 = shift_q_map_35;
      end
      6'b100100 : begin
        _zz_shift_q_6_8 = shift_q_map_36;
      end
      6'b100101 : begin
        _zz_shift_q_6_8 = shift_q_map_37;
      end
      6'b100110 : begin
        _zz_shift_q_6_8 = shift_q_map_38;
      end
      default : begin
        _zz_shift_q_6_8 = shift_q_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_i_7_9)
      6'b000000 : begin
        _zz_shift_i_7_8 = shift_i_map_0;
      end
      6'b000001 : begin
        _zz_shift_i_7_8 = shift_i_map_1;
      end
      6'b000010 : begin
        _zz_shift_i_7_8 = shift_i_map_2;
      end
      6'b000011 : begin
        _zz_shift_i_7_8 = shift_i_map_3;
      end
      6'b000100 : begin
        _zz_shift_i_7_8 = shift_i_map_4;
      end
      6'b000101 : begin
        _zz_shift_i_7_8 = shift_i_map_5;
      end
      6'b000110 : begin
        _zz_shift_i_7_8 = shift_i_map_6;
      end
      6'b000111 : begin
        _zz_shift_i_7_8 = shift_i_map_7;
      end
      6'b001000 : begin
        _zz_shift_i_7_8 = shift_i_map_8;
      end
      6'b001001 : begin
        _zz_shift_i_7_8 = shift_i_map_9;
      end
      6'b001010 : begin
        _zz_shift_i_7_8 = shift_i_map_10;
      end
      6'b001011 : begin
        _zz_shift_i_7_8 = shift_i_map_11;
      end
      6'b001100 : begin
        _zz_shift_i_7_8 = shift_i_map_12;
      end
      6'b001101 : begin
        _zz_shift_i_7_8 = shift_i_map_13;
      end
      6'b001110 : begin
        _zz_shift_i_7_8 = shift_i_map_14;
      end
      6'b001111 : begin
        _zz_shift_i_7_8 = shift_i_map_15;
      end
      6'b010000 : begin
        _zz_shift_i_7_8 = shift_i_map_16;
      end
      6'b010001 : begin
        _zz_shift_i_7_8 = shift_i_map_17;
      end
      6'b010010 : begin
        _zz_shift_i_7_8 = shift_i_map_18;
      end
      6'b010011 : begin
        _zz_shift_i_7_8 = shift_i_map_19;
      end
      6'b010100 : begin
        _zz_shift_i_7_8 = shift_i_map_20;
      end
      6'b010101 : begin
        _zz_shift_i_7_8 = shift_i_map_21;
      end
      6'b010110 : begin
        _zz_shift_i_7_8 = shift_i_map_22;
      end
      6'b010111 : begin
        _zz_shift_i_7_8 = shift_i_map_23;
      end
      6'b011000 : begin
        _zz_shift_i_7_8 = shift_i_map_24;
      end
      6'b011001 : begin
        _zz_shift_i_7_8 = shift_i_map_25;
      end
      6'b011010 : begin
        _zz_shift_i_7_8 = shift_i_map_26;
      end
      6'b011011 : begin
        _zz_shift_i_7_8 = shift_i_map_27;
      end
      6'b011100 : begin
        _zz_shift_i_7_8 = shift_i_map_28;
      end
      6'b011101 : begin
        _zz_shift_i_7_8 = shift_i_map_29;
      end
      6'b011110 : begin
        _zz_shift_i_7_8 = shift_i_map_30;
      end
      6'b011111 : begin
        _zz_shift_i_7_8 = shift_i_map_31;
      end
      6'b100000 : begin
        _zz_shift_i_7_8 = shift_i_map_32;
      end
      6'b100001 : begin
        _zz_shift_i_7_8 = shift_i_map_33;
      end
      6'b100010 : begin
        _zz_shift_i_7_8 = shift_i_map_34;
      end
      6'b100011 : begin
        _zz_shift_i_7_8 = shift_i_map_35;
      end
      6'b100100 : begin
        _zz_shift_i_7_8 = shift_i_map_36;
      end
      6'b100101 : begin
        _zz_shift_i_7_8 = shift_i_map_37;
      end
      6'b100110 : begin
        _zz_shift_i_7_8 = shift_i_map_38;
      end
      default : begin
        _zz_shift_i_7_8 = shift_i_map_39;
      end
    endcase
  end

  always @(*) begin
    case(_zz_shift_q_7_9)
      6'b000000 : begin
        _zz_shift_q_7_8 = shift_q_map_0;
      end
      6'b000001 : begin
        _zz_shift_q_7_8 = shift_q_map_1;
      end
      6'b000010 : begin
        _zz_shift_q_7_8 = shift_q_map_2;
      end
      6'b000011 : begin
        _zz_shift_q_7_8 = shift_q_map_3;
      end
      6'b000100 : begin
        _zz_shift_q_7_8 = shift_q_map_4;
      end
      6'b000101 : begin
        _zz_shift_q_7_8 = shift_q_map_5;
      end
      6'b000110 : begin
        _zz_shift_q_7_8 = shift_q_map_6;
      end
      6'b000111 : begin
        _zz_shift_q_7_8 = shift_q_map_7;
      end
      6'b001000 : begin
        _zz_shift_q_7_8 = shift_q_map_8;
      end
      6'b001001 : begin
        _zz_shift_q_7_8 = shift_q_map_9;
      end
      6'b001010 : begin
        _zz_shift_q_7_8 = shift_q_map_10;
      end
      6'b001011 : begin
        _zz_shift_q_7_8 = shift_q_map_11;
      end
      6'b001100 : begin
        _zz_shift_q_7_8 = shift_q_map_12;
      end
      6'b001101 : begin
        _zz_shift_q_7_8 = shift_q_map_13;
      end
      6'b001110 : begin
        _zz_shift_q_7_8 = shift_q_map_14;
      end
      6'b001111 : begin
        _zz_shift_q_7_8 = shift_q_map_15;
      end
      6'b010000 : begin
        _zz_shift_q_7_8 = shift_q_map_16;
      end
      6'b010001 : begin
        _zz_shift_q_7_8 = shift_q_map_17;
      end
      6'b010010 : begin
        _zz_shift_q_7_8 = shift_q_map_18;
      end
      6'b010011 : begin
        _zz_shift_q_7_8 = shift_q_map_19;
      end
      6'b010100 : begin
        _zz_shift_q_7_8 = shift_q_map_20;
      end
      6'b010101 : begin
        _zz_shift_q_7_8 = shift_q_map_21;
      end
      6'b010110 : begin
        _zz_shift_q_7_8 = shift_q_map_22;
      end
      6'b010111 : begin
        _zz_shift_q_7_8 = shift_q_map_23;
      end
      6'b011000 : begin
        _zz_shift_q_7_8 = shift_q_map_24;
      end
      6'b011001 : begin
        _zz_shift_q_7_8 = shift_q_map_25;
      end
      6'b011010 : begin
        _zz_shift_q_7_8 = shift_q_map_26;
      end
      6'b011011 : begin
        _zz_shift_q_7_8 = shift_q_map_27;
      end
      6'b011100 : begin
        _zz_shift_q_7_8 = shift_q_map_28;
      end
      6'b011101 : begin
        _zz_shift_q_7_8 = shift_q_map_29;
      end
      6'b011110 : begin
        _zz_shift_q_7_8 = shift_q_map_30;
      end
      6'b011111 : begin
        _zz_shift_q_7_8 = shift_q_map_31;
      end
      6'b100000 : begin
        _zz_shift_q_7_8 = shift_q_map_32;
      end
      6'b100001 : begin
        _zz_shift_q_7_8 = shift_q_map_33;
      end
      6'b100010 : begin
        _zz_shift_q_7_8 = shift_q_map_34;
      end
      6'b100011 : begin
        _zz_shift_q_7_8 = shift_q_map_35;
      end
      6'b100100 : begin
        _zz_shift_q_7_8 = shift_q_map_36;
      end
      6'b100101 : begin
        _zz_shift_q_7_8 = shift_q_map_37;
      end
      6'b100110 : begin
        _zz_shift_q_7_8 = shift_q_map_38;
      end
      default : begin
        _zz_shift_q_7_8 = shift_q_map_39;
      end
    endcase
  end

  assign _zz_1 = ({63'd0,1'b1} <<< w_addr);
  assign _zz_2 = ({63'd0,1'b1} <<< w_addr);
  assign base_sub_iqs_payload_0_cha_i = oAMUnspin_5_base_sub_iq_payload_cha_i;
  assign base_sub_iqs_payload_0_cha_q = oAMUnspin_5_base_sub_iq_payload_cha_q;
  assign base_sub_valid_vec_0 = oAMUnspin_5_base_sub_iq_valid;
  assign oAMUnspin_5_shift_i_0 = _zz_shift_i_0;
  assign oAMUnspin_5_shift_q_0 = _zz_shift_q_0;
  assign oAMUnspin_5_shift_i_1 = _zz_shift_i_1;
  assign oAMUnspin_5_shift_q_1 = _zz_shift_q_1;
  assign oAMUnspin_5_shift_i_2 = _zz_shift_i_2;
  assign oAMUnspin_5_shift_q_2 = _zz_shift_q_2;
  assign oAMUnspin_5_shift_i_3 = _zz_shift_i_3;
  assign oAMUnspin_5_shift_q_3 = _zz_shift_q_3;
  assign oAMUnspin_5_shift_i_4 = _zz_shift_i_4;
  assign oAMUnspin_5_shift_q_4 = _zz_shift_q_4;
  assign oAMUnspin_5_shift_i_5 = _zz_shift_i_5;
  assign oAMUnspin_5_shift_q_5 = _zz_shift_q_5;
  assign oAMUnspin_5_shift_i_6 = _zz_shift_i_6;
  assign oAMUnspin_5_shift_q_6 = _zz_shift_q_6;
  assign oAMUnspin_5_shift_i_7 = _zz_shift_i_7;
  assign oAMUnspin_5_shift_q_7 = _zz_shift_q_7;
  assign base_sub_iqs_payload_1_cha_i = oAMUnspin_6_base_sub_iq_payload_cha_i;
  assign base_sub_iqs_payload_1_cha_q = oAMUnspin_6_base_sub_iq_payload_cha_q;
  assign base_sub_valid_vec_1 = oAMUnspin_6_base_sub_iq_valid;
  assign oAMUnspin_6_shift_i_0 = _zz_shift_i_0_2;
  assign oAMUnspin_6_shift_q_0 = _zz_shift_q_0_2;
  assign oAMUnspin_6_shift_i_1 = _zz_shift_i_1_2;
  assign oAMUnspin_6_shift_q_1 = _zz_shift_q_1_2;
  assign oAMUnspin_6_shift_i_2 = _zz_shift_i_2_2;
  assign oAMUnspin_6_shift_q_2 = _zz_shift_q_2_2;
  assign oAMUnspin_6_shift_i_3 = _zz_shift_i_3_2;
  assign oAMUnspin_6_shift_q_3 = _zz_shift_q_3_2;
  assign oAMUnspin_6_shift_i_4 = _zz_shift_i_4_2;
  assign oAMUnspin_6_shift_q_4 = _zz_shift_q_4_2;
  assign oAMUnspin_6_shift_i_5 = _zz_shift_i_5_2;
  assign oAMUnspin_6_shift_q_5 = _zz_shift_q_5_2;
  assign oAMUnspin_6_shift_i_6 = _zz_shift_i_6_2;
  assign oAMUnspin_6_shift_q_6 = _zz_shift_q_6_2;
  assign oAMUnspin_6_shift_i_7 = _zz_shift_i_7_2;
  assign oAMUnspin_6_shift_q_7 = _zz_shift_q_7_2;
  assign base_sub_iqs_payload_2_cha_i = oAMUnspin_7_base_sub_iq_payload_cha_i;
  assign base_sub_iqs_payload_2_cha_q = oAMUnspin_7_base_sub_iq_payload_cha_q;
  assign base_sub_valid_vec_2 = oAMUnspin_7_base_sub_iq_valid;
  assign oAMUnspin_7_shift_i_0 = _zz_shift_i_0_4;
  assign oAMUnspin_7_shift_q_0 = _zz_shift_q_0_4;
  assign oAMUnspin_7_shift_i_1 = _zz_shift_i_1_4;
  assign oAMUnspin_7_shift_q_1 = _zz_shift_q_1_4;
  assign oAMUnspin_7_shift_i_2 = _zz_shift_i_2_4;
  assign oAMUnspin_7_shift_q_2 = _zz_shift_q_2_4;
  assign oAMUnspin_7_shift_i_3 = _zz_shift_i_3_4;
  assign oAMUnspin_7_shift_q_3 = _zz_shift_q_3_4;
  assign oAMUnspin_7_shift_i_4 = _zz_shift_i_4_4;
  assign oAMUnspin_7_shift_q_4 = _zz_shift_q_4_4;
  assign oAMUnspin_7_shift_i_5 = _zz_shift_i_5_4;
  assign oAMUnspin_7_shift_q_5 = _zz_shift_q_5_4;
  assign oAMUnspin_7_shift_i_6 = _zz_shift_i_6_4;
  assign oAMUnspin_7_shift_q_6 = _zz_shift_q_6_4;
  assign oAMUnspin_7_shift_i_7 = _zz_shift_i_7_4;
  assign oAMUnspin_7_shift_q_7 = _zz_shift_q_7_4;
  assign base_sub_iqs_payload_3_cha_i = oAMUnspin_8_base_sub_iq_payload_cha_i;
  assign base_sub_iqs_payload_3_cha_q = oAMUnspin_8_base_sub_iq_payload_cha_q;
  assign base_sub_valid_vec_3 = oAMUnspin_8_base_sub_iq_valid;
  assign oAMUnspin_8_shift_i_0 = _zz_shift_i_0_6;
  assign oAMUnspin_8_shift_q_0 = _zz_shift_q_0_6;
  assign oAMUnspin_8_shift_i_1 = _zz_shift_i_1_6;
  assign oAMUnspin_8_shift_q_1 = _zz_shift_q_1_6;
  assign oAMUnspin_8_shift_i_2 = _zz_shift_i_2_6;
  assign oAMUnspin_8_shift_q_2 = _zz_shift_q_2_6;
  assign oAMUnspin_8_shift_i_3 = _zz_shift_i_3_6;
  assign oAMUnspin_8_shift_q_3 = _zz_shift_q_3_6;
  assign oAMUnspin_8_shift_i_4 = _zz_shift_i_4_6;
  assign oAMUnspin_8_shift_q_4 = _zz_shift_q_4_6;
  assign oAMUnspin_8_shift_i_5 = _zz_shift_i_5_6;
  assign oAMUnspin_8_shift_q_5 = _zz_shift_q_5_6;
  assign oAMUnspin_8_shift_i_6 = _zz_shift_i_6_6;
  assign oAMUnspin_8_shift_q_6 = _zz_shift_q_6_6;
  assign oAMUnspin_8_shift_i_7 = _zz_shift_i_7_6;
  assign oAMUnspin_8_shift_q_7 = _zz_shift_q_7_6;
  assign base_sub_iqs_payload_4_cha_i = oAMUnspin_9_base_sub_iq_payload_cha_i;
  assign base_sub_iqs_payload_4_cha_q = oAMUnspin_9_base_sub_iq_payload_cha_q;
  assign base_sub_valid_vec_4 = oAMUnspin_9_base_sub_iq_valid;
  assign oAMUnspin_9_shift_i_0 = _zz_shift_i_0_8;
  assign oAMUnspin_9_shift_q_0 = _zz_shift_q_0_8;
  assign oAMUnspin_9_shift_i_1 = _zz_shift_i_1_8;
  assign oAMUnspin_9_shift_q_1 = _zz_shift_q_1_8;
  assign oAMUnspin_9_shift_i_2 = _zz_shift_i_2_8;
  assign oAMUnspin_9_shift_q_2 = _zz_shift_q_2_8;
  assign oAMUnspin_9_shift_i_3 = _zz_shift_i_3_8;
  assign oAMUnspin_9_shift_q_3 = _zz_shift_q_3_8;
  assign oAMUnspin_9_shift_i_4 = _zz_shift_i_4_8;
  assign oAMUnspin_9_shift_q_4 = _zz_shift_q_4_8;
  assign oAMUnspin_9_shift_i_5 = _zz_shift_i_5_8;
  assign oAMUnspin_9_shift_q_5 = _zz_shift_q_5_8;
  assign oAMUnspin_9_shift_i_6 = _zz_shift_i_6_8;
  assign oAMUnspin_9_shift_q_6 = _zz_shift_q_6_8;
  assign oAMUnspin_9_shift_i_7 = _zz_shift_i_7_8;
  assign oAMUnspin_9_shift_q_7 = _zz_shift_q_7_8;
  assign base_sub_iqs_valid = ((((base_sub_valid_vec_0 && base_sub_valid_vec_1) && base_sub_valid_vec_2) && base_sub_valid_vec_3) && base_sub_valid_vec_4);
  assign mod_iq_ready = (! w_en);
  always @(posedge clk) begin
    if(w_en) begin
      if(w_sel) begin
        if(_zz_1[0]) begin
          shift_i_map_0 <= w_data;
        end
        if(_zz_1[1]) begin
          shift_i_map_1 <= w_data;
        end
        if(_zz_1[2]) begin
          shift_i_map_2 <= w_data;
        end
        if(_zz_1[3]) begin
          shift_i_map_3 <= w_data;
        end
        if(_zz_1[4]) begin
          shift_i_map_4 <= w_data;
        end
        if(_zz_1[5]) begin
          shift_i_map_5 <= w_data;
        end
        if(_zz_1[6]) begin
          shift_i_map_6 <= w_data;
        end
        if(_zz_1[7]) begin
          shift_i_map_7 <= w_data;
        end
        if(_zz_1[8]) begin
          shift_i_map_8 <= w_data;
        end
        if(_zz_1[9]) begin
          shift_i_map_9 <= w_data;
        end
        if(_zz_1[10]) begin
          shift_i_map_10 <= w_data;
        end
        if(_zz_1[11]) begin
          shift_i_map_11 <= w_data;
        end
        if(_zz_1[12]) begin
          shift_i_map_12 <= w_data;
        end
        if(_zz_1[13]) begin
          shift_i_map_13 <= w_data;
        end
        if(_zz_1[14]) begin
          shift_i_map_14 <= w_data;
        end
        if(_zz_1[15]) begin
          shift_i_map_15 <= w_data;
        end
        if(_zz_1[16]) begin
          shift_i_map_16 <= w_data;
        end
        if(_zz_1[17]) begin
          shift_i_map_17 <= w_data;
        end
        if(_zz_1[18]) begin
          shift_i_map_18 <= w_data;
        end
        if(_zz_1[19]) begin
          shift_i_map_19 <= w_data;
        end
        if(_zz_1[20]) begin
          shift_i_map_20 <= w_data;
        end
        if(_zz_1[21]) begin
          shift_i_map_21 <= w_data;
        end
        if(_zz_1[22]) begin
          shift_i_map_22 <= w_data;
        end
        if(_zz_1[23]) begin
          shift_i_map_23 <= w_data;
        end
        if(_zz_1[24]) begin
          shift_i_map_24 <= w_data;
        end
        if(_zz_1[25]) begin
          shift_i_map_25 <= w_data;
        end
        if(_zz_1[26]) begin
          shift_i_map_26 <= w_data;
        end
        if(_zz_1[27]) begin
          shift_i_map_27 <= w_data;
        end
        if(_zz_1[28]) begin
          shift_i_map_28 <= w_data;
        end
        if(_zz_1[29]) begin
          shift_i_map_29 <= w_data;
        end
        if(_zz_1[30]) begin
          shift_i_map_30 <= w_data;
        end
        if(_zz_1[31]) begin
          shift_i_map_31 <= w_data;
        end
        if(_zz_1[32]) begin
          shift_i_map_32 <= w_data;
        end
        if(_zz_1[33]) begin
          shift_i_map_33 <= w_data;
        end
        if(_zz_1[34]) begin
          shift_i_map_34 <= w_data;
        end
        if(_zz_1[35]) begin
          shift_i_map_35 <= w_data;
        end
        if(_zz_1[36]) begin
          shift_i_map_36 <= w_data;
        end
        if(_zz_1[37]) begin
          shift_i_map_37 <= w_data;
        end
        if(_zz_1[38]) begin
          shift_i_map_38 <= w_data;
        end
        if(_zz_1[39]) begin
          shift_i_map_39 <= w_data;
        end
      end else begin
        if(_zz_2[0]) begin
          shift_q_map_0 <= w_data;
        end
        if(_zz_2[1]) begin
          shift_q_map_1 <= w_data;
        end
        if(_zz_2[2]) begin
          shift_q_map_2 <= w_data;
        end
        if(_zz_2[3]) begin
          shift_q_map_3 <= w_data;
        end
        if(_zz_2[4]) begin
          shift_q_map_4 <= w_data;
        end
        if(_zz_2[5]) begin
          shift_q_map_5 <= w_data;
        end
        if(_zz_2[6]) begin
          shift_q_map_6 <= w_data;
        end
        if(_zz_2[7]) begin
          shift_q_map_7 <= w_data;
        end
        if(_zz_2[8]) begin
          shift_q_map_8 <= w_data;
        end
        if(_zz_2[9]) begin
          shift_q_map_9 <= w_data;
        end
        if(_zz_2[10]) begin
          shift_q_map_10 <= w_data;
        end
        if(_zz_2[11]) begin
          shift_q_map_11 <= w_data;
        end
        if(_zz_2[12]) begin
          shift_q_map_12 <= w_data;
        end
        if(_zz_2[13]) begin
          shift_q_map_13 <= w_data;
        end
        if(_zz_2[14]) begin
          shift_q_map_14 <= w_data;
        end
        if(_zz_2[15]) begin
          shift_q_map_15 <= w_data;
        end
        if(_zz_2[16]) begin
          shift_q_map_16 <= w_data;
        end
        if(_zz_2[17]) begin
          shift_q_map_17 <= w_data;
        end
        if(_zz_2[18]) begin
          shift_q_map_18 <= w_data;
        end
        if(_zz_2[19]) begin
          shift_q_map_19 <= w_data;
        end
        if(_zz_2[20]) begin
          shift_q_map_20 <= w_data;
        end
        if(_zz_2[21]) begin
          shift_q_map_21 <= w_data;
        end
        if(_zz_2[22]) begin
          shift_q_map_22 <= w_data;
        end
        if(_zz_2[23]) begin
          shift_q_map_23 <= w_data;
        end
        if(_zz_2[24]) begin
          shift_q_map_24 <= w_data;
        end
        if(_zz_2[25]) begin
          shift_q_map_25 <= w_data;
        end
        if(_zz_2[26]) begin
          shift_q_map_26 <= w_data;
        end
        if(_zz_2[27]) begin
          shift_q_map_27 <= w_data;
        end
        if(_zz_2[28]) begin
          shift_q_map_28 <= w_data;
        end
        if(_zz_2[29]) begin
          shift_q_map_29 <= w_data;
        end
        if(_zz_2[30]) begin
          shift_q_map_30 <= w_data;
        end
        if(_zz_2[31]) begin
          shift_q_map_31 <= w_data;
        end
        if(_zz_2[32]) begin
          shift_q_map_32 <= w_data;
        end
        if(_zz_2[33]) begin
          shift_q_map_33 <= w_data;
        end
        if(_zz_2[34]) begin
          shift_q_map_34 <= w_data;
        end
        if(_zz_2[35]) begin
          shift_q_map_35 <= w_data;
        end
        if(_zz_2[36]) begin
          shift_q_map_36 <= w_data;
        end
        if(_zz_2[37]) begin
          shift_q_map_37 <= w_data;
        end
        if(_zz_2[38]) begin
          shift_q_map_38 <= w_data;
        end
        if(_zz_2[39]) begin
          shift_q_map_39 <= w_data;
        end
      end
    end
  end


endmodule

//OAMUnspin replaced by OAMUnspin

//OAMUnspin replaced by OAMUnspin

//OAMUnspin replaced by OAMUnspin

//OAMUnspin replaced by OAMUnspin

module OAMUnspin (
  input      [15:0]   shift_i_0,
  input      [15:0]   shift_i_1,
  input      [15:0]   shift_i_2,
  input      [15:0]   shift_i_3,
  input      [15:0]   shift_i_4,
  input      [15:0]   shift_i_5,
  input      [15:0]   shift_i_6,
  input      [15:0]   shift_i_7,
  input      [15:0]   shift_q_0,
  input      [15:0]   shift_q_1,
  input      [15:0]   shift_q_2,
  input      [15:0]   shift_q_3,
  input      [15:0]   shift_q_4,
  input      [15:0]   shift_q_5,
  input      [15:0]   shift_q_6,
  input      [15:0]   shift_q_7,
  input               mod_iq_valid,
  input      [15:0]   mod_iq_payload_cha_i,
  input      [15:0]   mod_iq_payload_cha_q,
  output              base_sub_iq_valid,
  output     [31:0]   base_sub_iq_payload_cha_i,
  output     [31:0]   base_sub_iq_payload_cha_q,
  input               clk,
  input               resetn
);
  wire       [31:0]   _zz_trans_i_vec_0;
  wire       [31:0]   _zz_trans_i_vec_0_1;
  wire       [31:0]   _zz_trans_q_vec_0;
  wire       [31:0]   _zz_trans_q_vec_0_1;
  wire       [31:0]   _zz_trans_i_vec_1;
  wire       [31:0]   _zz_trans_i_vec_1_1;
  wire       [31:0]   _zz_trans_q_vec_1;
  wire       [31:0]   _zz_trans_q_vec_1_1;
  wire       [31:0]   _zz_trans_i_vec_2;
  wire       [31:0]   _zz_trans_i_vec_2_1;
  wire       [31:0]   _zz_trans_q_vec_2;
  wire       [31:0]   _zz_trans_q_vec_2_1;
  wire       [31:0]   _zz_trans_i_vec_3;
  wire       [31:0]   _zz_trans_i_vec_3_1;
  wire       [31:0]   _zz_trans_q_vec_3;
  wire       [31:0]   _zz_trans_q_vec_3_1;
  wire       [31:0]   _zz_trans_i_vec_4;
  wire       [31:0]   _zz_trans_i_vec_4_1;
  wire       [31:0]   _zz_trans_q_vec_4;
  wire       [31:0]   _zz_trans_q_vec_4_1;
  wire       [31:0]   _zz_trans_i_vec_5;
  wire       [31:0]   _zz_trans_i_vec_5_1;
  wire       [31:0]   _zz_trans_q_vec_5;
  wire       [31:0]   _zz_trans_q_vec_5_1;
  wire       [31:0]   _zz_trans_i_vec_6;
  wire       [31:0]   _zz_trans_i_vec_6_1;
  wire       [31:0]   _zz_trans_q_vec_6;
  wire       [31:0]   _zz_trans_q_vec_6_1;
  wire       [31:0]   _zz_trans_i_vec_7;
  wire       [31:0]   _zz_trans_i_vec_7_1;
  wire       [31:0]   _zz_trans_q_vec_7;
  wire       [31:0]   _zz_trans_q_vec_7_1;
  wire       [30:0]   _zz__zz_base_sub_iq_payload_cha_i;
  wire       [31:0]   _zz__zz_base_sub_iq_payload_cha_i_1;
  wire       [30:0]   _zz__zz_base_sub_iq_payload_cha_i_1_1;
  wire       [31:0]   _zz__zz_base_sub_iq_payload_cha_i_1_2;
  wire       [30:0]   _zz__zz_base_sub_iq_payload_cha_i_2;
  wire       [31:0]   _zz__zz_base_sub_iq_payload_cha_i_2_1;
  wire       [30:0]   _zz__zz_base_sub_iq_payload_cha_i_3;
  wire       [31:0]   _zz__zz_base_sub_iq_payload_cha_i_3_1;
  wire       [30:0]   _zz__zz_base_sub_iq_payload_cha_i_4;
  wire       [31:0]   _zz__zz_base_sub_iq_payload_cha_i_4_1;
  wire       [30:0]   _zz__zz_base_sub_iq_payload_cha_i_5;
  wire       [31:0]   _zz__zz_base_sub_iq_payload_cha_i_5_1;
  wire       [30:0]   _zz__zz_base_sub_iq_payload_cha_i_6;
  wire       [31:0]   _zz__zz_base_sub_iq_payload_cha_i_6_1;
  wire       [30:0]   _zz__zz_base_sub_iq_payload_cha_q;
  wire       [31:0]   _zz__zz_base_sub_iq_payload_cha_q_1;
  wire       [30:0]   _zz__zz_base_sub_iq_payload_cha_q_1_1;
  wire       [31:0]   _zz__zz_base_sub_iq_payload_cha_q_1_2;
  wire       [30:0]   _zz__zz_base_sub_iq_payload_cha_q_2;
  wire       [31:0]   _zz__zz_base_sub_iq_payload_cha_q_2_1;
  wire       [30:0]   _zz__zz_base_sub_iq_payload_cha_q_3;
  wire       [31:0]   _zz__zz_base_sub_iq_payload_cha_q_3_1;
  wire       [30:0]   _zz__zz_base_sub_iq_payload_cha_q_4;
  wire       [31:0]   _zz__zz_base_sub_iq_payload_cha_q_4_1;
  wire       [30:0]   _zz__zz_base_sub_iq_payload_cha_q_5;
  wire       [31:0]   _zz__zz_base_sub_iq_payload_cha_q_5_1;
  wire       [30:0]   _zz__zz_base_sub_iq_payload_cha_q_6;
  wire       [31:0]   _zz__zz_base_sub_iq_payload_cha_q_6_1;
  reg        [15:0]   mod_iq_buf_cha_i;
  reg        [15:0]   mod_iq_buf_cha_q;
  reg                 mod_valid_buf;
  reg        [31:0]   trans_i_vec_0;
  reg        [31:0]   trans_i_vec_1;
  reg        [31:0]   trans_i_vec_2;
  reg        [31:0]   trans_i_vec_3;
  reg        [31:0]   trans_i_vec_4;
  reg        [31:0]   trans_i_vec_5;
  reg        [31:0]   trans_i_vec_6;
  reg        [31:0]   trans_i_vec_7;
  reg        [31:0]   trans_q_vec_0;
  reg        [31:0]   trans_q_vec_1;
  reg        [31:0]   trans_q_vec_2;
  reg        [31:0]   trans_q_vec_3;
  reg        [31:0]   trans_q_vec_4;
  reg        [31:0]   trans_q_vec_5;
  reg        [31:0]   trans_q_vec_6;
  reg        [31:0]   trans_q_vec_7;
  reg                 trans_valid;
  reg        [31:0]   _zz_base_sub_iq_payload_cha_i;
  reg        [31:0]   _zz_base_sub_iq_payload_cha_i_1;
  reg        [31:0]   _zz_base_sub_iq_payload_cha_i_2;
  reg        [31:0]   _zz_base_sub_iq_payload_cha_i_3;
  reg        [31:0]   _zz_base_sub_iq_payload_cha_i_4;
  reg        [31:0]   _zz_base_sub_iq_payload_cha_i_5;
  reg        [31:0]   _zz_base_sub_iq_payload_cha_i_6;
  reg        [31:0]   _zz_base_sub_iq_payload_cha_q;
  reg        [31:0]   _zz_base_sub_iq_payload_cha_q_1;
  reg        [31:0]   _zz_base_sub_iq_payload_cha_q_2;
  reg        [31:0]   _zz_base_sub_iq_payload_cha_q_3;
  reg        [31:0]   _zz_base_sub_iq_payload_cha_q_4;
  reg        [31:0]   _zz_base_sub_iq_payload_cha_q_5;
  reg        [31:0]   _zz_base_sub_iq_payload_cha_q_6;
  reg                 trans_valid_delay_1;
  reg                 trans_valid_delay_2;
  reg                 trans_valid_delay_3;

  assign _zz_trans_i_vec_0 = ($signed(mod_iq_buf_cha_i) * $signed(shift_i_0));
  assign _zz_trans_i_vec_0_1 = ($signed(mod_iq_buf_cha_q) * $signed(shift_q_0));
  assign _zz_trans_q_vec_0 = ($signed(mod_iq_buf_cha_i) * $signed(shift_q_0));
  assign _zz_trans_q_vec_0_1 = ($signed(mod_iq_buf_cha_q) * $signed(shift_i_0));
  assign _zz_trans_i_vec_1 = ($signed(mod_iq_buf_cha_i) * $signed(shift_i_1));
  assign _zz_trans_i_vec_1_1 = ($signed(mod_iq_buf_cha_q) * $signed(shift_q_1));
  assign _zz_trans_q_vec_1 = ($signed(mod_iq_buf_cha_i) * $signed(shift_q_1));
  assign _zz_trans_q_vec_1_1 = ($signed(mod_iq_buf_cha_q) * $signed(shift_i_1));
  assign _zz_trans_i_vec_2 = ($signed(mod_iq_buf_cha_i) * $signed(shift_i_2));
  assign _zz_trans_i_vec_2_1 = ($signed(mod_iq_buf_cha_q) * $signed(shift_q_2));
  assign _zz_trans_q_vec_2 = ($signed(mod_iq_buf_cha_i) * $signed(shift_q_2));
  assign _zz_trans_q_vec_2_1 = ($signed(mod_iq_buf_cha_q) * $signed(shift_i_2));
  assign _zz_trans_i_vec_3 = ($signed(mod_iq_buf_cha_i) * $signed(shift_i_3));
  assign _zz_trans_i_vec_3_1 = ($signed(mod_iq_buf_cha_q) * $signed(shift_q_3));
  assign _zz_trans_q_vec_3 = ($signed(mod_iq_buf_cha_i) * $signed(shift_q_3));
  assign _zz_trans_q_vec_3_1 = ($signed(mod_iq_buf_cha_q) * $signed(shift_i_3));
  assign _zz_trans_i_vec_4 = ($signed(mod_iq_buf_cha_i) * $signed(shift_i_4));
  assign _zz_trans_i_vec_4_1 = ($signed(mod_iq_buf_cha_q) * $signed(shift_q_4));
  assign _zz_trans_q_vec_4 = ($signed(mod_iq_buf_cha_i) * $signed(shift_q_4));
  assign _zz_trans_q_vec_4_1 = ($signed(mod_iq_buf_cha_q) * $signed(shift_i_4));
  assign _zz_trans_i_vec_5 = ($signed(mod_iq_buf_cha_i) * $signed(shift_i_5));
  assign _zz_trans_i_vec_5_1 = ($signed(mod_iq_buf_cha_q) * $signed(shift_q_5));
  assign _zz_trans_q_vec_5 = ($signed(mod_iq_buf_cha_i) * $signed(shift_q_5));
  assign _zz_trans_q_vec_5_1 = ($signed(mod_iq_buf_cha_q) * $signed(shift_i_5));
  assign _zz_trans_i_vec_6 = ($signed(mod_iq_buf_cha_i) * $signed(shift_i_6));
  assign _zz_trans_i_vec_6_1 = ($signed(mod_iq_buf_cha_q) * $signed(shift_q_6));
  assign _zz_trans_q_vec_6 = ($signed(mod_iq_buf_cha_i) * $signed(shift_q_6));
  assign _zz_trans_q_vec_6_1 = ($signed(mod_iq_buf_cha_q) * $signed(shift_i_6));
  assign _zz_trans_i_vec_7 = ($signed(mod_iq_buf_cha_i) * $signed(shift_i_7));
  assign _zz_trans_i_vec_7_1 = ($signed(mod_iq_buf_cha_q) * $signed(shift_q_7));
  assign _zz_trans_q_vec_7 = ($signed(mod_iq_buf_cha_i) * $signed(shift_q_7));
  assign _zz_trans_q_vec_7_1 = ($signed(mod_iq_buf_cha_q) * $signed(shift_i_7));
  assign _zz__zz_base_sub_iq_payload_cha_i = (_zz__zz_base_sub_iq_payload_cha_i_1 >>> 1);
  assign _zz__zz_base_sub_iq_payload_cha_i_1 = ($signed(trans_i_vec_0) + $signed(trans_i_vec_1));
  assign _zz__zz_base_sub_iq_payload_cha_i_1_1 = (_zz__zz_base_sub_iq_payload_cha_i_1_2 >>> 1);
  assign _zz__zz_base_sub_iq_payload_cha_i_1_2 = ($signed(trans_i_vec_2) + $signed(trans_i_vec_3));
  assign _zz__zz_base_sub_iq_payload_cha_i_2 = (_zz__zz_base_sub_iq_payload_cha_i_2_1 >>> 1);
  assign _zz__zz_base_sub_iq_payload_cha_i_2_1 = ($signed(trans_i_vec_4) + $signed(trans_i_vec_5));
  assign _zz__zz_base_sub_iq_payload_cha_i_3 = (_zz__zz_base_sub_iq_payload_cha_i_3_1 >>> 1);
  assign _zz__zz_base_sub_iq_payload_cha_i_3_1 = ($signed(trans_i_vec_6) + $signed(trans_i_vec_7));
  assign _zz__zz_base_sub_iq_payload_cha_i_4 = (_zz__zz_base_sub_iq_payload_cha_i_4_1 >>> 1);
  assign _zz__zz_base_sub_iq_payload_cha_i_4_1 = ($signed(_zz_base_sub_iq_payload_cha_i) + $signed(_zz_base_sub_iq_payload_cha_i_1));
  assign _zz__zz_base_sub_iq_payload_cha_i_5 = (_zz__zz_base_sub_iq_payload_cha_i_5_1 >>> 1);
  assign _zz__zz_base_sub_iq_payload_cha_i_5_1 = ($signed(_zz_base_sub_iq_payload_cha_i_2) + $signed(_zz_base_sub_iq_payload_cha_i_3));
  assign _zz__zz_base_sub_iq_payload_cha_i_6 = (_zz__zz_base_sub_iq_payload_cha_i_6_1 >>> 1);
  assign _zz__zz_base_sub_iq_payload_cha_i_6_1 = ($signed(_zz_base_sub_iq_payload_cha_i_4) + $signed(_zz_base_sub_iq_payload_cha_i_5));
  assign _zz__zz_base_sub_iq_payload_cha_q = (_zz__zz_base_sub_iq_payload_cha_q_1 >>> 1);
  assign _zz__zz_base_sub_iq_payload_cha_q_1 = ($signed(trans_q_vec_0) + $signed(trans_q_vec_1));
  assign _zz__zz_base_sub_iq_payload_cha_q_1_1 = (_zz__zz_base_sub_iq_payload_cha_q_1_2 >>> 1);
  assign _zz__zz_base_sub_iq_payload_cha_q_1_2 = ($signed(trans_q_vec_2) + $signed(trans_q_vec_3));
  assign _zz__zz_base_sub_iq_payload_cha_q_2 = (_zz__zz_base_sub_iq_payload_cha_q_2_1 >>> 1);
  assign _zz__zz_base_sub_iq_payload_cha_q_2_1 = ($signed(trans_q_vec_4) + $signed(trans_q_vec_5));
  assign _zz__zz_base_sub_iq_payload_cha_q_3 = (_zz__zz_base_sub_iq_payload_cha_q_3_1 >>> 1);
  assign _zz__zz_base_sub_iq_payload_cha_q_3_1 = ($signed(trans_q_vec_6) + $signed(trans_q_vec_7));
  assign _zz__zz_base_sub_iq_payload_cha_q_4 = (_zz__zz_base_sub_iq_payload_cha_q_4_1 >>> 1);
  assign _zz__zz_base_sub_iq_payload_cha_q_4_1 = ($signed(_zz_base_sub_iq_payload_cha_q) + $signed(_zz_base_sub_iq_payload_cha_q_1));
  assign _zz__zz_base_sub_iq_payload_cha_q_5 = (_zz__zz_base_sub_iq_payload_cha_q_5_1 >>> 1);
  assign _zz__zz_base_sub_iq_payload_cha_q_5_1 = ($signed(_zz_base_sub_iq_payload_cha_q_2) + $signed(_zz_base_sub_iq_payload_cha_q_3));
  assign _zz__zz_base_sub_iq_payload_cha_q_6 = (_zz__zz_base_sub_iq_payload_cha_q_6_1 >>> 1);
  assign _zz__zz_base_sub_iq_payload_cha_q_6_1 = ($signed(_zz_base_sub_iq_payload_cha_q_4) + $signed(_zz_base_sub_iq_payload_cha_q_5));
  assign base_sub_iq_payload_cha_i = _zz_base_sub_iq_payload_cha_i_6;
  assign base_sub_iq_payload_cha_q = _zz_base_sub_iq_payload_cha_q_6;
  assign base_sub_iq_valid = trans_valid_delay_3;
  always @(posedge clk) begin
    mod_iq_buf_cha_i <= mod_iq_payload_cha_i;
    mod_iq_buf_cha_q <= mod_iq_payload_cha_q;
    if(mod_valid_buf) begin
      trans_i_vec_0 <= ($signed(_zz_trans_i_vec_0) - $signed(_zz_trans_i_vec_0_1));
      trans_q_vec_0 <= ($signed(_zz_trans_q_vec_0) + $signed(_zz_trans_q_vec_0_1));
      trans_i_vec_1 <= ($signed(_zz_trans_i_vec_1) - $signed(_zz_trans_i_vec_1_1));
      trans_q_vec_1 <= ($signed(_zz_trans_q_vec_1) + $signed(_zz_trans_q_vec_1_1));
      trans_i_vec_2 <= ($signed(_zz_trans_i_vec_2) - $signed(_zz_trans_i_vec_2_1));
      trans_q_vec_2 <= ($signed(_zz_trans_q_vec_2) + $signed(_zz_trans_q_vec_2_1));
      trans_i_vec_3 <= ($signed(_zz_trans_i_vec_3) - $signed(_zz_trans_i_vec_3_1));
      trans_q_vec_3 <= ($signed(_zz_trans_q_vec_3) + $signed(_zz_trans_q_vec_3_1));
      trans_i_vec_4 <= ($signed(_zz_trans_i_vec_4) - $signed(_zz_trans_i_vec_4_1));
      trans_q_vec_4 <= ($signed(_zz_trans_q_vec_4) + $signed(_zz_trans_q_vec_4_1));
      trans_i_vec_5 <= ($signed(_zz_trans_i_vec_5) - $signed(_zz_trans_i_vec_5_1));
      trans_q_vec_5 <= ($signed(_zz_trans_q_vec_5) + $signed(_zz_trans_q_vec_5_1));
      trans_i_vec_6 <= ($signed(_zz_trans_i_vec_6) - $signed(_zz_trans_i_vec_6_1));
      trans_q_vec_6 <= ($signed(_zz_trans_q_vec_6) + $signed(_zz_trans_q_vec_6_1));
      trans_i_vec_7 <= ($signed(_zz_trans_i_vec_7) - $signed(_zz_trans_i_vec_7_1));
      trans_q_vec_7 <= ($signed(_zz_trans_q_vec_7) + $signed(_zz_trans_q_vec_7_1));
    end else begin
      trans_i_vec_0 <= 32'h0;
      trans_q_vec_0 <= 32'h0;
      trans_i_vec_1 <= 32'h0;
      trans_q_vec_1 <= 32'h0;
      trans_i_vec_2 <= 32'h0;
      trans_q_vec_2 <= 32'h0;
      trans_i_vec_3 <= 32'h0;
      trans_q_vec_3 <= 32'h0;
      trans_i_vec_4 <= 32'h0;
      trans_q_vec_4 <= 32'h0;
      trans_i_vec_5 <= 32'h0;
      trans_q_vec_5 <= 32'h0;
      trans_i_vec_6 <= 32'h0;
      trans_q_vec_6 <= 32'h0;
      trans_i_vec_7 <= 32'h0;
      trans_q_vec_7 <= 32'h0;
    end
    _zz_base_sub_iq_payload_cha_i <= {{1{_zz__zz_base_sub_iq_payload_cha_i[30]}}, _zz__zz_base_sub_iq_payload_cha_i};
    _zz_base_sub_iq_payload_cha_i_1 <= {{1{_zz__zz_base_sub_iq_payload_cha_i_1_1[30]}}, _zz__zz_base_sub_iq_payload_cha_i_1_1};
    _zz_base_sub_iq_payload_cha_i_2 <= {{1{_zz__zz_base_sub_iq_payload_cha_i_2[30]}}, _zz__zz_base_sub_iq_payload_cha_i_2};
    _zz_base_sub_iq_payload_cha_i_3 <= {{1{_zz__zz_base_sub_iq_payload_cha_i_3[30]}}, _zz__zz_base_sub_iq_payload_cha_i_3};
    _zz_base_sub_iq_payload_cha_i_4 <= {{1{_zz__zz_base_sub_iq_payload_cha_i_4[30]}}, _zz__zz_base_sub_iq_payload_cha_i_4};
    _zz_base_sub_iq_payload_cha_i_5 <= {{1{_zz__zz_base_sub_iq_payload_cha_i_5[30]}}, _zz__zz_base_sub_iq_payload_cha_i_5};
    _zz_base_sub_iq_payload_cha_i_6 <= {{1{_zz__zz_base_sub_iq_payload_cha_i_6[30]}}, _zz__zz_base_sub_iq_payload_cha_i_6};
    _zz_base_sub_iq_payload_cha_q <= {{1{_zz__zz_base_sub_iq_payload_cha_q[30]}}, _zz__zz_base_sub_iq_payload_cha_q};
    _zz_base_sub_iq_payload_cha_q_1 <= {{1{_zz__zz_base_sub_iq_payload_cha_q_1_1[30]}}, _zz__zz_base_sub_iq_payload_cha_q_1_1};
    _zz_base_sub_iq_payload_cha_q_2 <= {{1{_zz__zz_base_sub_iq_payload_cha_q_2[30]}}, _zz__zz_base_sub_iq_payload_cha_q_2};
    _zz_base_sub_iq_payload_cha_q_3 <= {{1{_zz__zz_base_sub_iq_payload_cha_q_3[30]}}, _zz__zz_base_sub_iq_payload_cha_q_3};
    _zz_base_sub_iq_payload_cha_q_4 <= {{1{_zz__zz_base_sub_iq_payload_cha_q_4[30]}}, _zz__zz_base_sub_iq_payload_cha_q_4};
    _zz_base_sub_iq_payload_cha_q_5 <= {{1{_zz__zz_base_sub_iq_payload_cha_q_5[30]}}, _zz__zz_base_sub_iq_payload_cha_q_5};
    _zz_base_sub_iq_payload_cha_q_6 <= {{1{_zz__zz_base_sub_iq_payload_cha_q_6[30]}}, _zz__zz_base_sub_iq_payload_cha_q_6};
    trans_valid_delay_1 <= trans_valid;
    trans_valid_delay_2 <= trans_valid_delay_1;
    trans_valid_delay_3 <= trans_valid_delay_2;
  end

  always @(posedge clk) begin
    if(!resetn) begin
      mod_valid_buf <= 1'b0;
      trans_valid <= 1'b0;
    end else begin
      mod_valid_buf <= mod_iq_valid;
      if(mod_valid_buf) begin
        trans_valid <= 1'b1;
      end else begin
        trans_valid <= 1'b0;
      end
    end
  end


endmodule
