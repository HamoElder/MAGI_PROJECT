// Generator : SpinalHDL v1.7.0    git head : eca519e78d4e6022e34911ec300a432ed9db8220
// Component : SystolicFIR
// Git hash  : fe8ed706a25b5cda33f96062d5bdc80425e016eb

`timescale 1ns/1ps

module SystolicFIR (
  input               raw_data_0_valid,
  input      [15:0]   raw_data_0_payload,
  input               raw_data_1_valid,
  input      [15:0]   raw_data_1_payload,
  input               raw_data_2_valid,
  input      [15:0]   raw_data_2_payload,
  input               raw_data_3_valid,
  input      [15:0]   raw_data_3_payload,
  output              filtered_data_0_valid,
  output     [31:0]   filtered_data_0_payload,
  output              filtered_data_1_valid,
  output     [31:0]   filtered_data_1_payload,
  output              filtered_data_2_valid,
  output     [31:0]   filtered_data_2_payload,
  output              filtered_data_3_valid,
  output     [31:0]   filtered_data_3_payload,
  input               clk,
  input               reset
);

  wire       [31:0]   systolicCore_116_input_data;
  wire       [31:0]   systolicCore_145_input_data;
  wire       [31:0]   systolicCore_174_input_data;
  wire       [31:0]   systolicCore_203_input_data;
  wire       [31:0]   systolicCore_116_next_input_data;
  wire       [31:0]   systolicCore_116_next_adder_data;
  wire                systolicCore_116_next_valid;
  wire       [31:0]   systolicCore_117_next_input_data;
  wire       [31:0]   systolicCore_117_next_adder_data;
  wire                systolicCore_117_next_valid;
  wire       [31:0]   systolicCore_118_next_input_data;
  wire       [31:0]   systolicCore_118_next_adder_data;
  wire                systolicCore_118_next_valid;
  wire       [31:0]   systolicCore_119_next_input_data;
  wire       [31:0]   systolicCore_119_next_adder_data;
  wire                systolicCore_119_next_valid;
  wire       [31:0]   systolicCore_120_next_input_data;
  wire       [31:0]   systolicCore_120_next_adder_data;
  wire                systolicCore_120_next_valid;
  wire       [31:0]   systolicCore_121_next_input_data;
  wire       [31:0]   systolicCore_121_next_adder_data;
  wire                systolicCore_121_next_valid;
  wire       [31:0]   systolicCore_122_next_input_data;
  wire       [31:0]   systolicCore_122_next_adder_data;
  wire                systolicCore_122_next_valid;
  wire       [31:0]   systolicCore_123_next_input_data;
  wire       [31:0]   systolicCore_123_next_adder_data;
  wire                systolicCore_123_next_valid;
  wire       [31:0]   systolicCore_124_next_input_data;
  wire       [31:0]   systolicCore_124_next_adder_data;
  wire                systolicCore_124_next_valid;
  wire       [31:0]   systolicCore_125_next_input_data;
  wire       [31:0]   systolicCore_125_next_adder_data;
  wire                systolicCore_125_next_valid;
  wire       [31:0]   systolicCore_126_next_input_data;
  wire       [31:0]   systolicCore_126_next_adder_data;
  wire                systolicCore_126_next_valid;
  wire       [31:0]   systolicCore_127_next_input_data;
  wire       [31:0]   systolicCore_127_next_adder_data;
  wire                systolicCore_127_next_valid;
  wire       [31:0]   systolicCore_128_next_input_data;
  wire       [31:0]   systolicCore_128_next_adder_data;
  wire                systolicCore_128_next_valid;
  wire       [31:0]   systolicCore_129_next_input_data;
  wire       [31:0]   systolicCore_129_next_adder_data;
  wire                systolicCore_129_next_valid;
  wire       [31:0]   systolicCore_130_next_input_data;
  wire       [31:0]   systolicCore_130_next_adder_data;
  wire                systolicCore_130_next_valid;
  wire       [31:0]   systolicCore_131_next_input_data;
  wire       [31:0]   systolicCore_131_next_adder_data;
  wire                systolicCore_131_next_valid;
  wire       [31:0]   systolicCore_132_next_input_data;
  wire       [31:0]   systolicCore_132_next_adder_data;
  wire                systolicCore_132_next_valid;
  wire       [31:0]   systolicCore_133_next_input_data;
  wire       [31:0]   systolicCore_133_next_adder_data;
  wire                systolicCore_133_next_valid;
  wire       [31:0]   systolicCore_134_next_input_data;
  wire       [31:0]   systolicCore_134_next_adder_data;
  wire                systolicCore_134_next_valid;
  wire       [31:0]   systolicCore_135_next_input_data;
  wire       [31:0]   systolicCore_135_next_adder_data;
  wire                systolicCore_135_next_valid;
  wire       [31:0]   systolicCore_136_next_input_data;
  wire       [31:0]   systolicCore_136_next_adder_data;
  wire                systolicCore_136_next_valid;
  wire       [31:0]   systolicCore_137_next_input_data;
  wire       [31:0]   systolicCore_137_next_adder_data;
  wire                systolicCore_137_next_valid;
  wire       [31:0]   systolicCore_138_next_input_data;
  wire       [31:0]   systolicCore_138_next_adder_data;
  wire                systolicCore_138_next_valid;
  wire       [31:0]   systolicCore_139_next_input_data;
  wire       [31:0]   systolicCore_139_next_adder_data;
  wire                systolicCore_139_next_valid;
  wire       [31:0]   systolicCore_140_next_input_data;
  wire       [31:0]   systolicCore_140_next_adder_data;
  wire                systolicCore_140_next_valid;
  wire       [31:0]   systolicCore_141_next_input_data;
  wire       [31:0]   systolicCore_141_next_adder_data;
  wire                systolicCore_141_next_valid;
  wire       [31:0]   systolicCore_142_next_input_data;
  wire       [31:0]   systolicCore_142_next_adder_data;
  wire                systolicCore_142_next_valid;
  wire       [31:0]   systolicCore_143_next_input_data;
  wire       [31:0]   systolicCore_143_next_adder_data;
  wire                systolicCore_143_next_valid;
  wire       [31:0]   systolicCore_144_next_input_data;
  wire       [31:0]   systolicCore_144_next_adder_data;
  wire                systolicCore_144_next_valid;
  wire       [31:0]   systolicCore_145_next_input_data;
  wire       [31:0]   systolicCore_145_next_adder_data;
  wire                systolicCore_145_next_valid;
  wire       [31:0]   systolicCore_146_next_input_data;
  wire       [31:0]   systolicCore_146_next_adder_data;
  wire                systolicCore_146_next_valid;
  wire       [31:0]   systolicCore_147_next_input_data;
  wire       [31:0]   systolicCore_147_next_adder_data;
  wire                systolicCore_147_next_valid;
  wire       [31:0]   systolicCore_148_next_input_data;
  wire       [31:0]   systolicCore_148_next_adder_data;
  wire                systolicCore_148_next_valid;
  wire       [31:0]   systolicCore_149_next_input_data;
  wire       [31:0]   systolicCore_149_next_adder_data;
  wire                systolicCore_149_next_valid;
  wire       [31:0]   systolicCore_150_next_input_data;
  wire       [31:0]   systolicCore_150_next_adder_data;
  wire                systolicCore_150_next_valid;
  wire       [31:0]   systolicCore_151_next_input_data;
  wire       [31:0]   systolicCore_151_next_adder_data;
  wire                systolicCore_151_next_valid;
  wire       [31:0]   systolicCore_152_next_input_data;
  wire       [31:0]   systolicCore_152_next_adder_data;
  wire                systolicCore_152_next_valid;
  wire       [31:0]   systolicCore_153_next_input_data;
  wire       [31:0]   systolicCore_153_next_adder_data;
  wire                systolicCore_153_next_valid;
  wire       [31:0]   systolicCore_154_next_input_data;
  wire       [31:0]   systolicCore_154_next_adder_data;
  wire                systolicCore_154_next_valid;
  wire       [31:0]   systolicCore_155_next_input_data;
  wire       [31:0]   systolicCore_155_next_adder_data;
  wire                systolicCore_155_next_valid;
  wire       [31:0]   systolicCore_156_next_input_data;
  wire       [31:0]   systolicCore_156_next_adder_data;
  wire                systolicCore_156_next_valid;
  wire       [31:0]   systolicCore_157_next_input_data;
  wire       [31:0]   systolicCore_157_next_adder_data;
  wire                systolicCore_157_next_valid;
  wire       [31:0]   systolicCore_158_next_input_data;
  wire       [31:0]   systolicCore_158_next_adder_data;
  wire                systolicCore_158_next_valid;
  wire       [31:0]   systolicCore_159_next_input_data;
  wire       [31:0]   systolicCore_159_next_adder_data;
  wire                systolicCore_159_next_valid;
  wire       [31:0]   systolicCore_160_next_input_data;
  wire       [31:0]   systolicCore_160_next_adder_data;
  wire                systolicCore_160_next_valid;
  wire       [31:0]   systolicCore_161_next_input_data;
  wire       [31:0]   systolicCore_161_next_adder_data;
  wire                systolicCore_161_next_valid;
  wire       [31:0]   systolicCore_162_next_input_data;
  wire       [31:0]   systolicCore_162_next_adder_data;
  wire                systolicCore_162_next_valid;
  wire       [31:0]   systolicCore_163_next_input_data;
  wire       [31:0]   systolicCore_163_next_adder_data;
  wire                systolicCore_163_next_valid;
  wire       [31:0]   systolicCore_164_next_input_data;
  wire       [31:0]   systolicCore_164_next_adder_data;
  wire                systolicCore_164_next_valid;
  wire       [31:0]   systolicCore_165_next_input_data;
  wire       [31:0]   systolicCore_165_next_adder_data;
  wire                systolicCore_165_next_valid;
  wire       [31:0]   systolicCore_166_next_input_data;
  wire       [31:0]   systolicCore_166_next_adder_data;
  wire                systolicCore_166_next_valid;
  wire       [31:0]   systolicCore_167_next_input_data;
  wire       [31:0]   systolicCore_167_next_adder_data;
  wire                systolicCore_167_next_valid;
  wire       [31:0]   systolicCore_168_next_input_data;
  wire       [31:0]   systolicCore_168_next_adder_data;
  wire                systolicCore_168_next_valid;
  wire       [31:0]   systolicCore_169_next_input_data;
  wire       [31:0]   systolicCore_169_next_adder_data;
  wire                systolicCore_169_next_valid;
  wire       [31:0]   systolicCore_170_next_input_data;
  wire       [31:0]   systolicCore_170_next_adder_data;
  wire                systolicCore_170_next_valid;
  wire       [31:0]   systolicCore_171_next_input_data;
  wire       [31:0]   systolicCore_171_next_adder_data;
  wire                systolicCore_171_next_valid;
  wire       [31:0]   systolicCore_172_next_input_data;
  wire       [31:0]   systolicCore_172_next_adder_data;
  wire                systolicCore_172_next_valid;
  wire       [31:0]   systolicCore_173_next_input_data;
  wire       [31:0]   systolicCore_173_next_adder_data;
  wire                systolicCore_173_next_valid;
  wire       [31:0]   systolicCore_174_next_input_data;
  wire       [31:0]   systolicCore_174_next_adder_data;
  wire                systolicCore_174_next_valid;
  wire       [31:0]   systolicCore_175_next_input_data;
  wire       [31:0]   systolicCore_175_next_adder_data;
  wire                systolicCore_175_next_valid;
  wire       [31:0]   systolicCore_176_next_input_data;
  wire       [31:0]   systolicCore_176_next_adder_data;
  wire                systolicCore_176_next_valid;
  wire       [31:0]   systolicCore_177_next_input_data;
  wire       [31:0]   systolicCore_177_next_adder_data;
  wire                systolicCore_177_next_valid;
  wire       [31:0]   systolicCore_178_next_input_data;
  wire       [31:0]   systolicCore_178_next_adder_data;
  wire                systolicCore_178_next_valid;
  wire       [31:0]   systolicCore_179_next_input_data;
  wire       [31:0]   systolicCore_179_next_adder_data;
  wire                systolicCore_179_next_valid;
  wire       [31:0]   systolicCore_180_next_input_data;
  wire       [31:0]   systolicCore_180_next_adder_data;
  wire                systolicCore_180_next_valid;
  wire       [31:0]   systolicCore_181_next_input_data;
  wire       [31:0]   systolicCore_181_next_adder_data;
  wire                systolicCore_181_next_valid;
  wire       [31:0]   systolicCore_182_next_input_data;
  wire       [31:0]   systolicCore_182_next_adder_data;
  wire                systolicCore_182_next_valid;
  wire       [31:0]   systolicCore_183_next_input_data;
  wire       [31:0]   systolicCore_183_next_adder_data;
  wire                systolicCore_183_next_valid;
  wire       [31:0]   systolicCore_184_next_input_data;
  wire       [31:0]   systolicCore_184_next_adder_data;
  wire                systolicCore_184_next_valid;
  wire       [31:0]   systolicCore_185_next_input_data;
  wire       [31:0]   systolicCore_185_next_adder_data;
  wire                systolicCore_185_next_valid;
  wire       [31:0]   systolicCore_186_next_input_data;
  wire       [31:0]   systolicCore_186_next_adder_data;
  wire                systolicCore_186_next_valid;
  wire       [31:0]   systolicCore_187_next_input_data;
  wire       [31:0]   systolicCore_187_next_adder_data;
  wire                systolicCore_187_next_valid;
  wire       [31:0]   systolicCore_188_next_input_data;
  wire       [31:0]   systolicCore_188_next_adder_data;
  wire                systolicCore_188_next_valid;
  wire       [31:0]   systolicCore_189_next_input_data;
  wire       [31:0]   systolicCore_189_next_adder_data;
  wire                systolicCore_189_next_valid;
  wire       [31:0]   systolicCore_190_next_input_data;
  wire       [31:0]   systolicCore_190_next_adder_data;
  wire                systolicCore_190_next_valid;
  wire       [31:0]   systolicCore_191_next_input_data;
  wire       [31:0]   systolicCore_191_next_adder_data;
  wire                systolicCore_191_next_valid;
  wire       [31:0]   systolicCore_192_next_input_data;
  wire       [31:0]   systolicCore_192_next_adder_data;
  wire                systolicCore_192_next_valid;
  wire       [31:0]   systolicCore_193_next_input_data;
  wire       [31:0]   systolicCore_193_next_adder_data;
  wire                systolicCore_193_next_valid;
  wire       [31:0]   systolicCore_194_next_input_data;
  wire       [31:0]   systolicCore_194_next_adder_data;
  wire                systolicCore_194_next_valid;
  wire       [31:0]   systolicCore_195_next_input_data;
  wire       [31:0]   systolicCore_195_next_adder_data;
  wire                systolicCore_195_next_valid;
  wire       [31:0]   systolicCore_196_next_input_data;
  wire       [31:0]   systolicCore_196_next_adder_data;
  wire                systolicCore_196_next_valid;
  wire       [31:0]   systolicCore_197_next_input_data;
  wire       [31:0]   systolicCore_197_next_adder_data;
  wire                systolicCore_197_next_valid;
  wire       [31:0]   systolicCore_198_next_input_data;
  wire       [31:0]   systolicCore_198_next_adder_data;
  wire                systolicCore_198_next_valid;
  wire       [31:0]   systolicCore_199_next_input_data;
  wire       [31:0]   systolicCore_199_next_adder_data;
  wire                systolicCore_199_next_valid;
  wire       [31:0]   systolicCore_200_next_input_data;
  wire       [31:0]   systolicCore_200_next_adder_data;
  wire                systolicCore_200_next_valid;
  wire       [31:0]   systolicCore_201_next_input_data;
  wire       [31:0]   systolicCore_201_next_adder_data;
  wire                systolicCore_201_next_valid;
  wire       [31:0]   systolicCore_202_next_input_data;
  wire       [31:0]   systolicCore_202_next_adder_data;
  wire                systolicCore_202_next_valid;
  wire       [31:0]   systolicCore_203_next_input_data;
  wire       [31:0]   systolicCore_203_next_adder_data;
  wire                systolicCore_203_next_valid;
  wire       [31:0]   systolicCore_204_next_input_data;
  wire       [31:0]   systolicCore_204_next_adder_data;
  wire                systolicCore_204_next_valid;
  wire       [31:0]   systolicCore_205_next_input_data;
  wire       [31:0]   systolicCore_205_next_adder_data;
  wire                systolicCore_205_next_valid;
  wire       [31:0]   systolicCore_206_next_input_data;
  wire       [31:0]   systolicCore_206_next_adder_data;
  wire                systolicCore_206_next_valid;
  wire       [31:0]   systolicCore_207_next_input_data;
  wire       [31:0]   systolicCore_207_next_adder_data;
  wire                systolicCore_207_next_valid;
  wire       [31:0]   systolicCore_208_next_input_data;
  wire       [31:0]   systolicCore_208_next_adder_data;
  wire                systolicCore_208_next_valid;
  wire       [31:0]   systolicCore_209_next_input_data;
  wire       [31:0]   systolicCore_209_next_adder_data;
  wire                systolicCore_209_next_valid;
  wire       [31:0]   systolicCore_210_next_input_data;
  wire       [31:0]   systolicCore_210_next_adder_data;
  wire                systolicCore_210_next_valid;
  wire       [31:0]   systolicCore_211_next_input_data;
  wire       [31:0]   systolicCore_211_next_adder_data;
  wire                systolicCore_211_next_valid;
  wire       [31:0]   systolicCore_212_next_input_data;
  wire       [31:0]   systolicCore_212_next_adder_data;
  wire                systolicCore_212_next_valid;
  wire       [31:0]   systolicCore_213_next_input_data;
  wire       [31:0]   systolicCore_213_next_adder_data;
  wire                systolicCore_213_next_valid;
  wire       [31:0]   systolicCore_214_next_input_data;
  wire       [31:0]   systolicCore_214_next_adder_data;
  wire                systolicCore_214_next_valid;
  wire       [31:0]   systolicCore_215_next_input_data;
  wire       [31:0]   systolicCore_215_next_adder_data;
  wire                systolicCore_215_next_valid;
  wire       [31:0]   systolicCore_216_next_input_data;
  wire       [31:0]   systolicCore_216_next_adder_data;
  wire                systolicCore_216_next_valid;
  wire       [31:0]   systolicCore_217_next_input_data;
  wire       [31:0]   systolicCore_217_next_adder_data;
  wire                systolicCore_217_next_valid;
  wire       [31:0]   systolicCore_218_next_input_data;
  wire       [31:0]   systolicCore_218_next_adder_data;
  wire                systolicCore_218_next_valid;
  wire       [31:0]   systolicCore_219_next_input_data;
  wire       [31:0]   systolicCore_219_next_adder_data;
  wire                systolicCore_219_next_valid;
  wire       [31:0]   systolicCore_220_next_input_data;
  wire       [31:0]   systolicCore_220_next_adder_data;
  wire                systolicCore_220_next_valid;
  wire       [31:0]   systolicCore_221_next_input_data;
  wire       [31:0]   systolicCore_221_next_adder_data;
  wire                systolicCore_221_next_valid;
  wire       [31:0]   systolicCore_222_next_input_data;
  wire       [31:0]   systolicCore_222_next_adder_data;
  wire                systolicCore_222_next_valid;
  wire       [31:0]   systolicCore_223_next_input_data;
  wire       [31:0]   systolicCore_223_next_adder_data;
  wire                systolicCore_223_next_valid;
  wire       [31:0]   systolicCore_224_next_input_data;
  wire       [31:0]   systolicCore_224_next_adder_data;
  wire                systolicCore_224_next_valid;
  wire       [31:0]   systolicCore_225_next_input_data;
  wire       [31:0]   systolicCore_225_next_adder_data;
  wire                systolicCore_225_next_valid;
  wire       [31:0]   systolicCore_226_next_input_data;
  wire       [31:0]   systolicCore_226_next_adder_data;
  wire                systolicCore_226_next_valid;
  wire       [31:0]   systolicCore_227_next_input_data;
  wire       [31:0]   systolicCore_227_next_adder_data;
  wire                systolicCore_227_next_valid;
  wire       [31:0]   systolicCore_228_next_input_data;
  wire       [31:0]   systolicCore_228_next_adder_data;
  wire                systolicCore_228_next_valid;
  wire       [31:0]   systolicCore_229_next_input_data;
  wire       [31:0]   systolicCore_229_next_adder_data;
  wire                systolicCore_229_next_valid;
  wire       [31:0]   systolicCore_230_next_input_data;
  wire       [31:0]   systolicCore_230_next_adder_data;
  wire                systolicCore_230_next_valid;
  wire       [31:0]   systolicCore_231_next_input_data;
  wire       [31:0]   systolicCore_231_next_adder_data;
  wire                systolicCore_231_next_valid;

  SystolicCore systolicCore_116 (
    .input_data      (systolicCore_116_input_data[31:0]     ), //i
    .coff_data       (6'h0                                  ), //i
    .adder_data      (32'h0                                 ), //i
    .valid           (raw_data_0_valid                      ), //i
    .next_input_data (systolicCore_116_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_116_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_116_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_117 (
    .input_data      (systolicCore_116_next_input_data[31:0]), //i
    .coff_data       (6'h0                                  ), //i
    .adder_data      (systolicCore_116_next_adder_data[31:0]), //i
    .valid           (systolicCore_116_next_valid           ), //i
    .next_input_data (systolicCore_117_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_117_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_117_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_118 (
    .input_data      (systolicCore_117_next_input_data[31:0]), //i
    .coff_data       (6'h0                                  ), //i
    .adder_data      (systolicCore_117_next_adder_data[31:0]), //i
    .valid           (systolicCore_117_next_valid           ), //i
    .next_input_data (systolicCore_118_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_118_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_118_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_119 (
    .input_data      (systolicCore_118_next_input_data[31:0]), //i
    .coff_data       (6'h01                                 ), //i
    .adder_data      (systolicCore_118_next_adder_data[31:0]), //i
    .valid           (systolicCore_118_next_valid           ), //i
    .next_input_data (systolicCore_119_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_119_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_119_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_120 (
    .input_data      (systolicCore_119_next_input_data[31:0]), //i
    .coff_data       (6'h01                                 ), //i
    .adder_data      (systolicCore_119_next_adder_data[31:0]), //i
    .valid           (systolicCore_119_next_valid           ), //i
    .next_input_data (systolicCore_120_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_120_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_120_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_121 (
    .input_data      (systolicCore_120_next_input_data[31:0]), //i
    .coff_data       (6'h03                                 ), //i
    .adder_data      (systolicCore_120_next_adder_data[31:0]), //i
    .valid           (systolicCore_120_next_valid           ), //i
    .next_input_data (systolicCore_121_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_121_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_121_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_122 (
    .input_data      (systolicCore_121_next_input_data[31:0]), //i
    .coff_data       (6'h05                                 ), //i
    .adder_data      (systolicCore_121_next_adder_data[31:0]), //i
    .valid           (systolicCore_121_next_valid           ), //i
    .next_input_data (systolicCore_122_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_122_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_122_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_123 (
    .input_data      (systolicCore_122_next_input_data[31:0]), //i
    .coff_data       (6'h07                                 ), //i
    .adder_data      (systolicCore_122_next_adder_data[31:0]), //i
    .valid           (systolicCore_122_next_valid           ), //i
    .next_input_data (systolicCore_123_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_123_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_123_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_124 (
    .input_data      (systolicCore_123_next_input_data[31:0]), //i
    .coff_data       (6'h0a                                 ), //i
    .adder_data      (systolicCore_123_next_adder_data[31:0]), //i
    .valid           (systolicCore_123_next_valid           ), //i
    .next_input_data (systolicCore_124_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_124_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_124_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_125 (
    .input_data      (systolicCore_124_next_input_data[31:0]), //i
    .coff_data       (6'h0d                                 ), //i
    .adder_data      (systolicCore_124_next_adder_data[31:0]), //i
    .valid           (systolicCore_124_next_valid           ), //i
    .next_input_data (systolicCore_125_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_125_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_125_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_126 (
    .input_data      (systolicCore_125_next_input_data[31:0]), //i
    .coff_data       (6'h10                                 ), //i
    .adder_data      (systolicCore_125_next_adder_data[31:0]), //i
    .valid           (systolicCore_125_next_valid           ), //i
    .next_input_data (systolicCore_126_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_126_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_126_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_127 (
    .input_data      (systolicCore_126_next_input_data[31:0]), //i
    .coff_data       (6'h13                                 ), //i
    .adder_data      (systolicCore_126_next_adder_data[31:0]), //i
    .valid           (systolicCore_126_next_valid           ), //i
    .next_input_data (systolicCore_127_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_127_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_127_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_128 (
    .input_data      (systolicCore_127_next_input_data[31:0]), //i
    .coff_data       (6'h15                                 ), //i
    .adder_data      (systolicCore_127_next_adder_data[31:0]), //i
    .valid           (systolicCore_127_next_valid           ), //i
    .next_input_data (systolicCore_128_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_128_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_128_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_129 (
    .input_data      (systolicCore_128_next_input_data[31:0]), //i
    .coff_data       (6'h17                                 ), //i
    .adder_data      (systolicCore_128_next_adder_data[31:0]), //i
    .valid           (systolicCore_128_next_valid           ), //i
    .next_input_data (systolicCore_129_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_129_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_129_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_130 (
    .input_data      (systolicCore_129_next_input_data[31:0]), //i
    .coff_data       (6'h17                                 ), //i
    .adder_data      (systolicCore_129_next_adder_data[31:0]), //i
    .valid           (systolicCore_129_next_valid           ), //i
    .next_input_data (systolicCore_130_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_130_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_130_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_131 (
    .input_data      (systolicCore_130_next_input_data[31:0]), //i
    .coff_data       (6'h17                                 ), //i
    .adder_data      (systolicCore_130_next_adder_data[31:0]), //i
    .valid           (systolicCore_130_next_valid           ), //i
    .next_input_data (systolicCore_131_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_131_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_131_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_132 (
    .input_data      (systolicCore_131_next_input_data[31:0]), //i
    .coff_data       (6'h15                                 ), //i
    .adder_data      (systolicCore_131_next_adder_data[31:0]), //i
    .valid           (systolicCore_131_next_valid           ), //i
    .next_input_data (systolicCore_132_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_132_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_132_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_133 (
    .input_data      (systolicCore_132_next_input_data[31:0]), //i
    .coff_data       (6'h13                                 ), //i
    .adder_data      (systolicCore_132_next_adder_data[31:0]), //i
    .valid           (systolicCore_132_next_valid           ), //i
    .next_input_data (systolicCore_133_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_133_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_133_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_134 (
    .input_data      (systolicCore_133_next_input_data[31:0]), //i
    .coff_data       (6'h10                                 ), //i
    .adder_data      (systolicCore_133_next_adder_data[31:0]), //i
    .valid           (systolicCore_133_next_valid           ), //i
    .next_input_data (systolicCore_134_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_134_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_134_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_135 (
    .input_data      (systolicCore_134_next_input_data[31:0]), //i
    .coff_data       (6'h0d                                 ), //i
    .adder_data      (systolicCore_134_next_adder_data[31:0]), //i
    .valid           (systolicCore_134_next_valid           ), //i
    .next_input_data (systolicCore_135_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_135_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_135_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_136 (
    .input_data      (systolicCore_135_next_input_data[31:0]), //i
    .coff_data       (6'h0a                                 ), //i
    .adder_data      (systolicCore_135_next_adder_data[31:0]), //i
    .valid           (systolicCore_135_next_valid           ), //i
    .next_input_data (systolicCore_136_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_136_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_136_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_137 (
    .input_data      (systolicCore_136_next_input_data[31:0]), //i
    .coff_data       (6'h07                                 ), //i
    .adder_data      (systolicCore_136_next_adder_data[31:0]), //i
    .valid           (systolicCore_136_next_valid           ), //i
    .next_input_data (systolicCore_137_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_137_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_137_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_138 (
    .input_data      (systolicCore_137_next_input_data[31:0]), //i
    .coff_data       (6'h05                                 ), //i
    .adder_data      (systolicCore_137_next_adder_data[31:0]), //i
    .valid           (systolicCore_137_next_valid           ), //i
    .next_input_data (systolicCore_138_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_138_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_138_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_139 (
    .input_data      (systolicCore_138_next_input_data[31:0]), //i
    .coff_data       (6'h03                                 ), //i
    .adder_data      (systolicCore_138_next_adder_data[31:0]), //i
    .valid           (systolicCore_138_next_valid           ), //i
    .next_input_data (systolicCore_139_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_139_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_139_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_140 (
    .input_data      (systolicCore_139_next_input_data[31:0]), //i
    .coff_data       (6'h01                                 ), //i
    .adder_data      (systolicCore_139_next_adder_data[31:0]), //i
    .valid           (systolicCore_139_next_valid           ), //i
    .next_input_data (systolicCore_140_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_140_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_140_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_141 (
    .input_data      (systolicCore_140_next_input_data[31:0]), //i
    .coff_data       (6'h01                                 ), //i
    .adder_data      (systolicCore_140_next_adder_data[31:0]), //i
    .valid           (systolicCore_140_next_valid           ), //i
    .next_input_data (systolicCore_141_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_141_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_141_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_142 (
    .input_data      (systolicCore_141_next_input_data[31:0]), //i
    .coff_data       (6'h0                                  ), //i
    .adder_data      (systolicCore_141_next_adder_data[31:0]), //i
    .valid           (systolicCore_141_next_valid           ), //i
    .next_input_data (systolicCore_142_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_142_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_142_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_143 (
    .input_data      (systolicCore_142_next_input_data[31:0]), //i
    .coff_data       (6'h0                                  ), //i
    .adder_data      (systolicCore_142_next_adder_data[31:0]), //i
    .valid           (systolicCore_142_next_valid           ), //i
    .next_input_data (systolicCore_143_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_143_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_143_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_144 (
    .input_data      (systolicCore_143_next_input_data[31:0]), //i
    .coff_data       (6'h0                                  ), //i
    .adder_data      (systolicCore_143_next_adder_data[31:0]), //i
    .valid           (systolicCore_143_next_valid           ), //i
    .next_input_data (systolicCore_144_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_144_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_144_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_145 (
    .input_data      (systolicCore_145_input_data[31:0]     ), //i
    .coff_data       (6'h0                                  ), //i
    .adder_data      (32'h0                                 ), //i
    .valid           (raw_data_1_valid                      ), //i
    .next_input_data (systolicCore_145_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_145_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_145_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_146 (
    .input_data      (systolicCore_145_next_input_data[31:0]), //i
    .coff_data       (6'h0                                  ), //i
    .adder_data      (systolicCore_145_next_adder_data[31:0]), //i
    .valid           (systolicCore_145_next_valid           ), //i
    .next_input_data (systolicCore_146_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_146_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_146_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_147 (
    .input_data      (systolicCore_146_next_input_data[31:0]), //i
    .coff_data       (6'h0                                  ), //i
    .adder_data      (systolicCore_146_next_adder_data[31:0]), //i
    .valid           (systolicCore_146_next_valid           ), //i
    .next_input_data (systolicCore_147_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_147_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_147_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_148 (
    .input_data      (systolicCore_147_next_input_data[31:0]), //i
    .coff_data       (6'h01                                 ), //i
    .adder_data      (systolicCore_147_next_adder_data[31:0]), //i
    .valid           (systolicCore_147_next_valid           ), //i
    .next_input_data (systolicCore_148_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_148_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_148_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_149 (
    .input_data      (systolicCore_148_next_input_data[31:0]), //i
    .coff_data       (6'h01                                 ), //i
    .adder_data      (systolicCore_148_next_adder_data[31:0]), //i
    .valid           (systolicCore_148_next_valid           ), //i
    .next_input_data (systolicCore_149_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_149_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_149_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_150 (
    .input_data      (systolicCore_149_next_input_data[31:0]), //i
    .coff_data       (6'h03                                 ), //i
    .adder_data      (systolicCore_149_next_adder_data[31:0]), //i
    .valid           (systolicCore_149_next_valid           ), //i
    .next_input_data (systolicCore_150_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_150_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_150_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_151 (
    .input_data      (systolicCore_150_next_input_data[31:0]), //i
    .coff_data       (6'h05                                 ), //i
    .adder_data      (systolicCore_150_next_adder_data[31:0]), //i
    .valid           (systolicCore_150_next_valid           ), //i
    .next_input_data (systolicCore_151_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_151_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_151_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_152 (
    .input_data      (systolicCore_151_next_input_data[31:0]), //i
    .coff_data       (6'h07                                 ), //i
    .adder_data      (systolicCore_151_next_adder_data[31:0]), //i
    .valid           (systolicCore_151_next_valid           ), //i
    .next_input_data (systolicCore_152_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_152_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_152_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_153 (
    .input_data      (systolicCore_152_next_input_data[31:0]), //i
    .coff_data       (6'h0a                                 ), //i
    .adder_data      (systolicCore_152_next_adder_data[31:0]), //i
    .valid           (systolicCore_152_next_valid           ), //i
    .next_input_data (systolicCore_153_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_153_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_153_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_154 (
    .input_data      (systolicCore_153_next_input_data[31:0]), //i
    .coff_data       (6'h0d                                 ), //i
    .adder_data      (systolicCore_153_next_adder_data[31:0]), //i
    .valid           (systolicCore_153_next_valid           ), //i
    .next_input_data (systolicCore_154_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_154_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_154_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_155 (
    .input_data      (systolicCore_154_next_input_data[31:0]), //i
    .coff_data       (6'h10                                 ), //i
    .adder_data      (systolicCore_154_next_adder_data[31:0]), //i
    .valid           (systolicCore_154_next_valid           ), //i
    .next_input_data (systolicCore_155_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_155_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_155_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_156 (
    .input_data      (systolicCore_155_next_input_data[31:0]), //i
    .coff_data       (6'h13                                 ), //i
    .adder_data      (systolicCore_155_next_adder_data[31:0]), //i
    .valid           (systolicCore_155_next_valid           ), //i
    .next_input_data (systolicCore_156_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_156_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_156_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_157 (
    .input_data      (systolicCore_156_next_input_data[31:0]), //i
    .coff_data       (6'h15                                 ), //i
    .adder_data      (systolicCore_156_next_adder_data[31:0]), //i
    .valid           (systolicCore_156_next_valid           ), //i
    .next_input_data (systolicCore_157_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_157_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_157_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_158 (
    .input_data      (systolicCore_157_next_input_data[31:0]), //i
    .coff_data       (6'h17                                 ), //i
    .adder_data      (systolicCore_157_next_adder_data[31:0]), //i
    .valid           (systolicCore_157_next_valid           ), //i
    .next_input_data (systolicCore_158_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_158_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_158_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_159 (
    .input_data      (systolicCore_158_next_input_data[31:0]), //i
    .coff_data       (6'h17                                 ), //i
    .adder_data      (systolicCore_158_next_adder_data[31:0]), //i
    .valid           (systolicCore_158_next_valid           ), //i
    .next_input_data (systolicCore_159_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_159_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_159_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_160 (
    .input_data      (systolicCore_159_next_input_data[31:0]), //i
    .coff_data       (6'h17                                 ), //i
    .adder_data      (systolicCore_159_next_adder_data[31:0]), //i
    .valid           (systolicCore_159_next_valid           ), //i
    .next_input_data (systolicCore_160_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_160_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_160_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_161 (
    .input_data      (systolicCore_160_next_input_data[31:0]), //i
    .coff_data       (6'h15                                 ), //i
    .adder_data      (systolicCore_160_next_adder_data[31:0]), //i
    .valid           (systolicCore_160_next_valid           ), //i
    .next_input_data (systolicCore_161_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_161_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_161_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_162 (
    .input_data      (systolicCore_161_next_input_data[31:0]), //i
    .coff_data       (6'h13                                 ), //i
    .adder_data      (systolicCore_161_next_adder_data[31:0]), //i
    .valid           (systolicCore_161_next_valid           ), //i
    .next_input_data (systolicCore_162_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_162_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_162_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_163 (
    .input_data      (systolicCore_162_next_input_data[31:0]), //i
    .coff_data       (6'h10                                 ), //i
    .adder_data      (systolicCore_162_next_adder_data[31:0]), //i
    .valid           (systolicCore_162_next_valid           ), //i
    .next_input_data (systolicCore_163_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_163_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_163_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_164 (
    .input_data      (systolicCore_163_next_input_data[31:0]), //i
    .coff_data       (6'h0d                                 ), //i
    .adder_data      (systolicCore_163_next_adder_data[31:0]), //i
    .valid           (systolicCore_163_next_valid           ), //i
    .next_input_data (systolicCore_164_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_164_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_164_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_165 (
    .input_data      (systolicCore_164_next_input_data[31:0]), //i
    .coff_data       (6'h0a                                 ), //i
    .adder_data      (systolicCore_164_next_adder_data[31:0]), //i
    .valid           (systolicCore_164_next_valid           ), //i
    .next_input_data (systolicCore_165_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_165_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_165_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_166 (
    .input_data      (systolicCore_165_next_input_data[31:0]), //i
    .coff_data       (6'h07                                 ), //i
    .adder_data      (systolicCore_165_next_adder_data[31:0]), //i
    .valid           (systolicCore_165_next_valid           ), //i
    .next_input_data (systolicCore_166_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_166_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_166_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_167 (
    .input_data      (systolicCore_166_next_input_data[31:0]), //i
    .coff_data       (6'h05                                 ), //i
    .adder_data      (systolicCore_166_next_adder_data[31:0]), //i
    .valid           (systolicCore_166_next_valid           ), //i
    .next_input_data (systolicCore_167_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_167_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_167_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_168 (
    .input_data      (systolicCore_167_next_input_data[31:0]), //i
    .coff_data       (6'h03                                 ), //i
    .adder_data      (systolicCore_167_next_adder_data[31:0]), //i
    .valid           (systolicCore_167_next_valid           ), //i
    .next_input_data (systolicCore_168_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_168_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_168_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_169 (
    .input_data      (systolicCore_168_next_input_data[31:0]), //i
    .coff_data       (6'h01                                 ), //i
    .adder_data      (systolicCore_168_next_adder_data[31:0]), //i
    .valid           (systolicCore_168_next_valid           ), //i
    .next_input_data (systolicCore_169_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_169_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_169_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_170 (
    .input_data      (systolicCore_169_next_input_data[31:0]), //i
    .coff_data       (6'h01                                 ), //i
    .adder_data      (systolicCore_169_next_adder_data[31:0]), //i
    .valid           (systolicCore_169_next_valid           ), //i
    .next_input_data (systolicCore_170_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_170_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_170_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_171 (
    .input_data      (systolicCore_170_next_input_data[31:0]), //i
    .coff_data       (6'h0                                  ), //i
    .adder_data      (systolicCore_170_next_adder_data[31:0]), //i
    .valid           (systolicCore_170_next_valid           ), //i
    .next_input_data (systolicCore_171_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_171_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_171_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_172 (
    .input_data      (systolicCore_171_next_input_data[31:0]), //i
    .coff_data       (6'h0                                  ), //i
    .adder_data      (systolicCore_171_next_adder_data[31:0]), //i
    .valid           (systolicCore_171_next_valid           ), //i
    .next_input_data (systolicCore_172_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_172_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_172_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_173 (
    .input_data      (systolicCore_172_next_input_data[31:0]), //i
    .coff_data       (6'h0                                  ), //i
    .adder_data      (systolicCore_172_next_adder_data[31:0]), //i
    .valid           (systolicCore_172_next_valid           ), //i
    .next_input_data (systolicCore_173_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_173_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_173_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_174 (
    .input_data      (systolicCore_174_input_data[31:0]     ), //i
    .coff_data       (6'h0                                  ), //i
    .adder_data      (32'h0                                 ), //i
    .valid           (raw_data_2_valid                      ), //i
    .next_input_data (systolicCore_174_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_174_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_174_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_175 (
    .input_data      (systolicCore_174_next_input_data[31:0]), //i
    .coff_data       (6'h0                                  ), //i
    .adder_data      (systolicCore_174_next_adder_data[31:0]), //i
    .valid           (systolicCore_174_next_valid           ), //i
    .next_input_data (systolicCore_175_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_175_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_175_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_176 (
    .input_data      (systolicCore_175_next_input_data[31:0]), //i
    .coff_data       (6'h0                                  ), //i
    .adder_data      (systolicCore_175_next_adder_data[31:0]), //i
    .valid           (systolicCore_175_next_valid           ), //i
    .next_input_data (systolicCore_176_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_176_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_176_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_177 (
    .input_data      (systolicCore_176_next_input_data[31:0]), //i
    .coff_data       (6'h01                                 ), //i
    .adder_data      (systolicCore_176_next_adder_data[31:0]), //i
    .valid           (systolicCore_176_next_valid           ), //i
    .next_input_data (systolicCore_177_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_177_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_177_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_178 (
    .input_data      (systolicCore_177_next_input_data[31:0]), //i
    .coff_data       (6'h01                                 ), //i
    .adder_data      (systolicCore_177_next_adder_data[31:0]), //i
    .valid           (systolicCore_177_next_valid           ), //i
    .next_input_data (systolicCore_178_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_178_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_178_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_179 (
    .input_data      (systolicCore_178_next_input_data[31:0]), //i
    .coff_data       (6'h03                                 ), //i
    .adder_data      (systolicCore_178_next_adder_data[31:0]), //i
    .valid           (systolicCore_178_next_valid           ), //i
    .next_input_data (systolicCore_179_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_179_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_179_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_180 (
    .input_data      (systolicCore_179_next_input_data[31:0]), //i
    .coff_data       (6'h05                                 ), //i
    .adder_data      (systolicCore_179_next_adder_data[31:0]), //i
    .valid           (systolicCore_179_next_valid           ), //i
    .next_input_data (systolicCore_180_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_180_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_180_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_181 (
    .input_data      (systolicCore_180_next_input_data[31:0]), //i
    .coff_data       (6'h07                                 ), //i
    .adder_data      (systolicCore_180_next_adder_data[31:0]), //i
    .valid           (systolicCore_180_next_valid           ), //i
    .next_input_data (systolicCore_181_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_181_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_181_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_182 (
    .input_data      (systolicCore_181_next_input_data[31:0]), //i
    .coff_data       (6'h0a                                 ), //i
    .adder_data      (systolicCore_181_next_adder_data[31:0]), //i
    .valid           (systolicCore_181_next_valid           ), //i
    .next_input_data (systolicCore_182_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_182_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_182_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_183 (
    .input_data      (systolicCore_182_next_input_data[31:0]), //i
    .coff_data       (6'h0d                                 ), //i
    .adder_data      (systolicCore_182_next_adder_data[31:0]), //i
    .valid           (systolicCore_182_next_valid           ), //i
    .next_input_data (systolicCore_183_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_183_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_183_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_184 (
    .input_data      (systolicCore_183_next_input_data[31:0]), //i
    .coff_data       (6'h10                                 ), //i
    .adder_data      (systolicCore_183_next_adder_data[31:0]), //i
    .valid           (systolicCore_183_next_valid           ), //i
    .next_input_data (systolicCore_184_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_184_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_184_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_185 (
    .input_data      (systolicCore_184_next_input_data[31:0]), //i
    .coff_data       (6'h13                                 ), //i
    .adder_data      (systolicCore_184_next_adder_data[31:0]), //i
    .valid           (systolicCore_184_next_valid           ), //i
    .next_input_data (systolicCore_185_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_185_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_185_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_186 (
    .input_data      (systolicCore_185_next_input_data[31:0]), //i
    .coff_data       (6'h15                                 ), //i
    .adder_data      (systolicCore_185_next_adder_data[31:0]), //i
    .valid           (systolicCore_185_next_valid           ), //i
    .next_input_data (systolicCore_186_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_186_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_186_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_187 (
    .input_data      (systolicCore_186_next_input_data[31:0]), //i
    .coff_data       (6'h17                                 ), //i
    .adder_data      (systolicCore_186_next_adder_data[31:0]), //i
    .valid           (systolicCore_186_next_valid           ), //i
    .next_input_data (systolicCore_187_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_187_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_187_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_188 (
    .input_data      (systolicCore_187_next_input_data[31:0]), //i
    .coff_data       (6'h17                                 ), //i
    .adder_data      (systolicCore_187_next_adder_data[31:0]), //i
    .valid           (systolicCore_187_next_valid           ), //i
    .next_input_data (systolicCore_188_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_188_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_188_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_189 (
    .input_data      (systolicCore_188_next_input_data[31:0]), //i
    .coff_data       (6'h17                                 ), //i
    .adder_data      (systolicCore_188_next_adder_data[31:0]), //i
    .valid           (systolicCore_188_next_valid           ), //i
    .next_input_data (systolicCore_189_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_189_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_189_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_190 (
    .input_data      (systolicCore_189_next_input_data[31:0]), //i
    .coff_data       (6'h15                                 ), //i
    .adder_data      (systolicCore_189_next_adder_data[31:0]), //i
    .valid           (systolicCore_189_next_valid           ), //i
    .next_input_data (systolicCore_190_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_190_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_190_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_191 (
    .input_data      (systolicCore_190_next_input_data[31:0]), //i
    .coff_data       (6'h13                                 ), //i
    .adder_data      (systolicCore_190_next_adder_data[31:0]), //i
    .valid           (systolicCore_190_next_valid           ), //i
    .next_input_data (systolicCore_191_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_191_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_191_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_192 (
    .input_data      (systolicCore_191_next_input_data[31:0]), //i
    .coff_data       (6'h10                                 ), //i
    .adder_data      (systolicCore_191_next_adder_data[31:0]), //i
    .valid           (systolicCore_191_next_valid           ), //i
    .next_input_data (systolicCore_192_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_192_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_192_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_193 (
    .input_data      (systolicCore_192_next_input_data[31:0]), //i
    .coff_data       (6'h0d                                 ), //i
    .adder_data      (systolicCore_192_next_adder_data[31:0]), //i
    .valid           (systolicCore_192_next_valid           ), //i
    .next_input_data (systolicCore_193_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_193_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_193_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_194 (
    .input_data      (systolicCore_193_next_input_data[31:0]), //i
    .coff_data       (6'h0a                                 ), //i
    .adder_data      (systolicCore_193_next_adder_data[31:0]), //i
    .valid           (systolicCore_193_next_valid           ), //i
    .next_input_data (systolicCore_194_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_194_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_194_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_195 (
    .input_data      (systolicCore_194_next_input_data[31:0]), //i
    .coff_data       (6'h07                                 ), //i
    .adder_data      (systolicCore_194_next_adder_data[31:0]), //i
    .valid           (systolicCore_194_next_valid           ), //i
    .next_input_data (systolicCore_195_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_195_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_195_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_196 (
    .input_data      (systolicCore_195_next_input_data[31:0]), //i
    .coff_data       (6'h05                                 ), //i
    .adder_data      (systolicCore_195_next_adder_data[31:0]), //i
    .valid           (systolicCore_195_next_valid           ), //i
    .next_input_data (systolicCore_196_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_196_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_196_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_197 (
    .input_data      (systolicCore_196_next_input_data[31:0]), //i
    .coff_data       (6'h03                                 ), //i
    .adder_data      (systolicCore_196_next_adder_data[31:0]), //i
    .valid           (systolicCore_196_next_valid           ), //i
    .next_input_data (systolicCore_197_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_197_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_197_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_198 (
    .input_data      (systolicCore_197_next_input_data[31:0]), //i
    .coff_data       (6'h01                                 ), //i
    .adder_data      (systolicCore_197_next_adder_data[31:0]), //i
    .valid           (systolicCore_197_next_valid           ), //i
    .next_input_data (systolicCore_198_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_198_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_198_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_199 (
    .input_data      (systolicCore_198_next_input_data[31:0]), //i
    .coff_data       (6'h01                                 ), //i
    .adder_data      (systolicCore_198_next_adder_data[31:0]), //i
    .valid           (systolicCore_198_next_valid           ), //i
    .next_input_data (systolicCore_199_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_199_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_199_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_200 (
    .input_data      (systolicCore_199_next_input_data[31:0]), //i
    .coff_data       (6'h0                                  ), //i
    .adder_data      (systolicCore_199_next_adder_data[31:0]), //i
    .valid           (systolicCore_199_next_valid           ), //i
    .next_input_data (systolicCore_200_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_200_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_200_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_201 (
    .input_data      (systolicCore_200_next_input_data[31:0]), //i
    .coff_data       (6'h0                                  ), //i
    .adder_data      (systolicCore_200_next_adder_data[31:0]), //i
    .valid           (systolicCore_200_next_valid           ), //i
    .next_input_data (systolicCore_201_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_201_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_201_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_202 (
    .input_data      (systolicCore_201_next_input_data[31:0]), //i
    .coff_data       (6'h0                                  ), //i
    .adder_data      (systolicCore_201_next_adder_data[31:0]), //i
    .valid           (systolicCore_201_next_valid           ), //i
    .next_input_data (systolicCore_202_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_202_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_202_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_203 (
    .input_data      (systolicCore_203_input_data[31:0]     ), //i
    .coff_data       (6'h0                                  ), //i
    .adder_data      (32'h0                                 ), //i
    .valid           (raw_data_3_valid                      ), //i
    .next_input_data (systolicCore_203_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_203_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_203_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_204 (
    .input_data      (systolicCore_203_next_input_data[31:0]), //i
    .coff_data       (6'h0                                  ), //i
    .adder_data      (systolicCore_203_next_adder_data[31:0]), //i
    .valid           (systolicCore_203_next_valid           ), //i
    .next_input_data (systolicCore_204_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_204_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_204_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_205 (
    .input_data      (systolicCore_204_next_input_data[31:0]), //i
    .coff_data       (6'h0                                  ), //i
    .adder_data      (systolicCore_204_next_adder_data[31:0]), //i
    .valid           (systolicCore_204_next_valid           ), //i
    .next_input_data (systolicCore_205_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_205_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_205_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_206 (
    .input_data      (systolicCore_205_next_input_data[31:0]), //i
    .coff_data       (6'h01                                 ), //i
    .adder_data      (systolicCore_205_next_adder_data[31:0]), //i
    .valid           (systolicCore_205_next_valid           ), //i
    .next_input_data (systolicCore_206_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_206_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_206_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_207 (
    .input_data      (systolicCore_206_next_input_data[31:0]), //i
    .coff_data       (6'h01                                 ), //i
    .adder_data      (systolicCore_206_next_adder_data[31:0]), //i
    .valid           (systolicCore_206_next_valid           ), //i
    .next_input_data (systolicCore_207_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_207_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_207_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_208 (
    .input_data      (systolicCore_207_next_input_data[31:0]), //i
    .coff_data       (6'h03                                 ), //i
    .adder_data      (systolicCore_207_next_adder_data[31:0]), //i
    .valid           (systolicCore_207_next_valid           ), //i
    .next_input_data (systolicCore_208_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_208_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_208_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_209 (
    .input_data      (systolicCore_208_next_input_data[31:0]), //i
    .coff_data       (6'h05                                 ), //i
    .adder_data      (systolicCore_208_next_adder_data[31:0]), //i
    .valid           (systolicCore_208_next_valid           ), //i
    .next_input_data (systolicCore_209_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_209_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_209_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_210 (
    .input_data      (systolicCore_209_next_input_data[31:0]), //i
    .coff_data       (6'h07                                 ), //i
    .adder_data      (systolicCore_209_next_adder_data[31:0]), //i
    .valid           (systolicCore_209_next_valid           ), //i
    .next_input_data (systolicCore_210_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_210_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_210_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_211 (
    .input_data      (systolicCore_210_next_input_data[31:0]), //i
    .coff_data       (6'h0a                                 ), //i
    .adder_data      (systolicCore_210_next_adder_data[31:0]), //i
    .valid           (systolicCore_210_next_valid           ), //i
    .next_input_data (systolicCore_211_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_211_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_211_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_212 (
    .input_data      (systolicCore_211_next_input_data[31:0]), //i
    .coff_data       (6'h0d                                 ), //i
    .adder_data      (systolicCore_211_next_adder_data[31:0]), //i
    .valid           (systolicCore_211_next_valid           ), //i
    .next_input_data (systolicCore_212_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_212_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_212_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_213 (
    .input_data      (systolicCore_212_next_input_data[31:0]), //i
    .coff_data       (6'h10                                 ), //i
    .adder_data      (systolicCore_212_next_adder_data[31:0]), //i
    .valid           (systolicCore_212_next_valid           ), //i
    .next_input_data (systolicCore_213_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_213_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_213_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_214 (
    .input_data      (systolicCore_213_next_input_data[31:0]), //i
    .coff_data       (6'h13                                 ), //i
    .adder_data      (systolicCore_213_next_adder_data[31:0]), //i
    .valid           (systolicCore_213_next_valid           ), //i
    .next_input_data (systolicCore_214_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_214_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_214_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_215 (
    .input_data      (systolicCore_214_next_input_data[31:0]), //i
    .coff_data       (6'h15                                 ), //i
    .adder_data      (systolicCore_214_next_adder_data[31:0]), //i
    .valid           (systolicCore_214_next_valid           ), //i
    .next_input_data (systolicCore_215_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_215_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_215_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_216 (
    .input_data      (systolicCore_215_next_input_data[31:0]), //i
    .coff_data       (6'h17                                 ), //i
    .adder_data      (systolicCore_215_next_adder_data[31:0]), //i
    .valid           (systolicCore_215_next_valid           ), //i
    .next_input_data (systolicCore_216_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_216_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_216_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_217 (
    .input_data      (systolicCore_216_next_input_data[31:0]), //i
    .coff_data       (6'h17                                 ), //i
    .adder_data      (systolicCore_216_next_adder_data[31:0]), //i
    .valid           (systolicCore_216_next_valid           ), //i
    .next_input_data (systolicCore_217_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_217_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_217_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_218 (
    .input_data      (systolicCore_217_next_input_data[31:0]), //i
    .coff_data       (6'h17                                 ), //i
    .adder_data      (systolicCore_217_next_adder_data[31:0]), //i
    .valid           (systolicCore_217_next_valid           ), //i
    .next_input_data (systolicCore_218_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_218_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_218_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_219 (
    .input_data      (systolicCore_218_next_input_data[31:0]), //i
    .coff_data       (6'h15                                 ), //i
    .adder_data      (systolicCore_218_next_adder_data[31:0]), //i
    .valid           (systolicCore_218_next_valid           ), //i
    .next_input_data (systolicCore_219_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_219_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_219_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_220 (
    .input_data      (systolicCore_219_next_input_data[31:0]), //i
    .coff_data       (6'h13                                 ), //i
    .adder_data      (systolicCore_219_next_adder_data[31:0]), //i
    .valid           (systolicCore_219_next_valid           ), //i
    .next_input_data (systolicCore_220_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_220_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_220_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_221 (
    .input_data      (systolicCore_220_next_input_data[31:0]), //i
    .coff_data       (6'h10                                 ), //i
    .adder_data      (systolicCore_220_next_adder_data[31:0]), //i
    .valid           (systolicCore_220_next_valid           ), //i
    .next_input_data (systolicCore_221_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_221_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_221_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_222 (
    .input_data      (systolicCore_221_next_input_data[31:0]), //i
    .coff_data       (6'h0d                                 ), //i
    .adder_data      (systolicCore_221_next_adder_data[31:0]), //i
    .valid           (systolicCore_221_next_valid           ), //i
    .next_input_data (systolicCore_222_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_222_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_222_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_223 (
    .input_data      (systolicCore_222_next_input_data[31:0]), //i
    .coff_data       (6'h0a                                 ), //i
    .adder_data      (systolicCore_222_next_adder_data[31:0]), //i
    .valid           (systolicCore_222_next_valid           ), //i
    .next_input_data (systolicCore_223_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_223_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_223_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_224 (
    .input_data      (systolicCore_223_next_input_data[31:0]), //i
    .coff_data       (6'h07                                 ), //i
    .adder_data      (systolicCore_223_next_adder_data[31:0]), //i
    .valid           (systolicCore_223_next_valid           ), //i
    .next_input_data (systolicCore_224_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_224_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_224_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_225 (
    .input_data      (systolicCore_224_next_input_data[31:0]), //i
    .coff_data       (6'h05                                 ), //i
    .adder_data      (systolicCore_224_next_adder_data[31:0]), //i
    .valid           (systolicCore_224_next_valid           ), //i
    .next_input_data (systolicCore_225_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_225_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_225_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_226 (
    .input_data      (systolicCore_225_next_input_data[31:0]), //i
    .coff_data       (6'h03                                 ), //i
    .adder_data      (systolicCore_225_next_adder_data[31:0]), //i
    .valid           (systolicCore_225_next_valid           ), //i
    .next_input_data (systolicCore_226_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_226_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_226_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_227 (
    .input_data      (systolicCore_226_next_input_data[31:0]), //i
    .coff_data       (6'h01                                 ), //i
    .adder_data      (systolicCore_226_next_adder_data[31:0]), //i
    .valid           (systolicCore_226_next_valid           ), //i
    .next_input_data (systolicCore_227_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_227_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_227_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_228 (
    .input_data      (systolicCore_227_next_input_data[31:0]), //i
    .coff_data       (6'h01                                 ), //i
    .adder_data      (systolicCore_227_next_adder_data[31:0]), //i
    .valid           (systolicCore_227_next_valid           ), //i
    .next_input_data (systolicCore_228_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_228_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_228_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_229 (
    .input_data      (systolicCore_228_next_input_data[31:0]), //i
    .coff_data       (6'h0                                  ), //i
    .adder_data      (systolicCore_228_next_adder_data[31:0]), //i
    .valid           (systolicCore_228_next_valid           ), //i
    .next_input_data (systolicCore_229_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_229_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_229_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_230 (
    .input_data      (systolicCore_229_next_input_data[31:0]), //i
    .coff_data       (6'h0                                  ), //i
    .adder_data      (systolicCore_229_next_adder_data[31:0]), //i
    .valid           (systolicCore_229_next_valid           ), //i
    .next_input_data (systolicCore_230_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_230_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_230_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  SystolicCore systolicCore_231 (
    .input_data      (systolicCore_230_next_input_data[31:0]), //i
    .coff_data       (6'h0                                  ), //i
    .adder_data      (systolicCore_230_next_adder_data[31:0]), //i
    .valid           (systolicCore_230_next_valid           ), //i
    .next_input_data (systolicCore_231_next_input_data[31:0]), //o
    .next_adder_data (systolicCore_231_next_adder_data[31:0]), //o
    .next_valid      (systolicCore_231_next_valid           ), //o
    .clk             (clk                                   ), //i
    .reset           (reset                                 )  //i
  );
  assign systolicCore_116_input_data = {{16{raw_data_0_payload[15]}}, raw_data_0_payload};
  assign filtered_data_0_payload = systolicCore_144_next_adder_data;
  assign filtered_data_0_valid = systolicCore_144_next_valid;
  assign systolicCore_145_input_data = {{16{raw_data_1_payload[15]}}, raw_data_1_payload};
  assign filtered_data_1_payload = systolicCore_173_next_adder_data;
  assign filtered_data_1_valid = systolicCore_173_next_valid;
  assign systolicCore_174_input_data = {{16{raw_data_2_payload[15]}}, raw_data_2_payload};
  assign filtered_data_2_payload = systolicCore_202_next_adder_data;
  assign filtered_data_2_valid = systolicCore_202_next_valid;
  assign systolicCore_203_input_data = {{16{raw_data_3_payload[15]}}, raw_data_3_payload};
  assign filtered_data_3_payload = systolicCore_231_next_adder_data;
  assign filtered_data_3_valid = systolicCore_231_next_valid;

endmodule

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

//SystolicCore replaced by SystolicCore

module SystolicCore (
  input      [31:0]   input_data,
  input      [5:0]    coff_data,
  input      [31:0]   adder_data,
  input               valid,
  output     [31:0]   next_input_data,
  output     [31:0]   next_adder_data,
  output              next_valid,
  input               clk,
  input               reset
);

  wire       [31:0]   shiftRegister_116_output_1;
  wire       [37:0]   _zz_next_adder;
  reg        [37:0]   mult;
  reg        [37:0]   next_adder;
  reg                 valid_regNext;

  assign _zz_next_adder = {{6{adder_data[31]}}, adder_data};
  ShiftRegister shiftRegister_116 (
    .input_1  (input_data[31:0]                ), //i
    .output_1 (shiftRegister_116_output_1[31:0]), //o
    .enable   (valid                           ), //i
    .clk      (clk                             ), //i
    .reset    (reset                           )  //i
  );
  assign next_valid = valid_regNext;
  assign next_input_data = shiftRegister_116_output_1;
  assign next_adder_data = next_adder[31:0];
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      mult <= 38'h0;
      next_adder <= 38'h0;
      valid_regNext <= 1'b0;
    end else begin
      if(valid) begin
        mult <= ($signed(coff_data) * $signed(shiftRegister_116_output_1));
      end
      if(valid) begin
        next_adder <= ($signed(mult) + $signed(_zz_next_adder));
      end
      valid_regNext <= valid;
    end
  end


endmodule

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

module ShiftRegister (
  input      [31:0]   input_1,
  output     [31:0]   output_1,
  input               enable,
  input               clk,
  input               reset
);

  reg        [31:0]   shift_reg_0;
  reg        [31:0]   shift_reg_1;

  assign output_1 = shift_reg_1;
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      shift_reg_0 <= 32'h0;
      shift_reg_1 <= 32'h0;
    end else begin
      if(enable) begin
        shift_reg_0 <= input_1;
        shift_reg_1 <= shift_reg_0;
      end
    end
  end


endmodule
