// Generator : SpinalHDL v1.6.0    git head : 73c8d8e2b86b45646e9d0b2e729291f2b65e6be3
// Component : R2MDC
// Git hash  : e3a5df1ea47c224930d57c25c9d0d9fb2bdff661



module R2MDC (
  input               mode,
  input               raw_data_valid,
  output              raw_data_ready,
  input      [23:0]   raw_data_payload_re,
  input      [23:0]   raw_data_payload_im,
  output              result_valid,
  output              result_payload_last,
  output     [23:0]   result_payload_fragment_re,
  output     [23:0]   result_payload_fragment_im,
  input               clk,
  input               reset
);
  wire       [23:0]   r2Butterfly_10_wn_re;
  wire       [23:0]   r2Butterfly_10_wn_im;
  wire                r2Switch_10_sel;
  wire       [23:0]   r2Butterfly_11_wn_re;
  wire       [23:0]   r2Butterfly_11_wn_im;
  wire                r2Switch_11_sel;
  wire       [23:0]   r2Butterfly_12_wn_re;
  wire       [23:0]   r2Butterfly_12_wn_im;
  wire                r2Switch_12_sel;
  wire       [23:0]   r2Butterfly_13_wn_re;
  wire       [23:0]   r2Butterfly_13_wn_im;
  wire                r2Switch_13_sel;
  wire       [23:0]   r2Butterfly_14_wn_re;
  wire       [23:0]   r2Butterfly_14_wn_im;
  wire                r2Switch_14_sel;
  wire       [23:0]   r2Butterfly_15_wn_re;
  wire       [23:0]   r2Butterfly_15_wn_im;
  wire                r2Switch_15_sel;
  wire       [23:0]   r2Butterfly_16_wn_re;
  wire       [23:0]   r2Butterfly_16_wn_im;
  wire                r2Switch_16_sel;
  wire       [23:0]   r2Butterfly_17_wn_re;
  wire       [23:0]   r2Butterfly_17_wn_im;
  wire                r2Switch_17_sel;
  wire       [23:0]   r2Butterfly_18_wn_re;
  wire       [23:0]   r2Butterfly_18_wn_im;
  wire                r2Switch_18_sel;
  wire       [23:0]   r2Butterfly_19_wn_re;
  wire       [23:0]   r2Butterfly_19_wn_im;
  wire                r2Switch_19_sel;
  wire                reorder_1_unsorted_valid;
  reg        [47:0]   _zz__zz_1_port0;
  reg        [47:0]   _zz__zz_2_port0;
  reg        [47:0]   _zz__zz_3_port0;
  reg        [47:0]   _zz__zz_4_port0;
  reg        [47:0]   _zz__zz_5_port0;
  reg        [47:0]   _zz__zz_6_port0;
  reg        [47:0]   _zz__zz_7_port0;
  reg        [47:0]   _zz__zz_8_port0;
  reg        [47:0]   _zz__zz_9_port0;
  reg        [47:0]   _zz__zz_10_port0;
  wire       [23:0]   shiftRegisterNE_20_output_re;
  wire       [23:0]   shiftRegisterNE_20_output_im;
  wire       [23:0]   r2Butterfly_10_out1_re;
  wire       [23:0]   r2Butterfly_10_out1_im;
  wire       [23:0]   r2Butterfly_10_out2_re;
  wire       [23:0]   r2Butterfly_10_out2_im;
  wire       [23:0]   shiftRegisterNE_21_output_re;
  wire       [23:0]   shiftRegisterNE_21_output_im;
  wire       [23:0]   r2Switch_10_out1_re;
  wire       [23:0]   r2Switch_10_out1_im;
  wire       [23:0]   r2Switch_10_out2_re;
  wire       [23:0]   r2Switch_10_out2_im;
  wire       [23:0]   shiftRegisterNE_22_output_re;
  wire       [23:0]   shiftRegisterNE_22_output_im;
  wire       [23:0]   r2Butterfly_11_out1_re;
  wire       [23:0]   r2Butterfly_11_out1_im;
  wire       [23:0]   r2Butterfly_11_out2_re;
  wire       [23:0]   r2Butterfly_11_out2_im;
  wire       [23:0]   shiftRegisterNE_23_output_re;
  wire       [23:0]   shiftRegisterNE_23_output_im;
  wire       [23:0]   r2Switch_11_out1_re;
  wire       [23:0]   r2Switch_11_out1_im;
  wire       [23:0]   r2Switch_11_out2_re;
  wire       [23:0]   r2Switch_11_out2_im;
  wire       [23:0]   shiftRegisterNE_24_output_re;
  wire       [23:0]   shiftRegisterNE_24_output_im;
  wire       [23:0]   r2Butterfly_12_out1_re;
  wire       [23:0]   r2Butterfly_12_out1_im;
  wire       [23:0]   r2Butterfly_12_out2_re;
  wire       [23:0]   r2Butterfly_12_out2_im;
  wire       [23:0]   shiftRegisterNE_25_output_re;
  wire       [23:0]   shiftRegisterNE_25_output_im;
  wire       [23:0]   r2Switch_12_out1_re;
  wire       [23:0]   r2Switch_12_out1_im;
  wire       [23:0]   r2Switch_12_out2_re;
  wire       [23:0]   r2Switch_12_out2_im;
  wire       [23:0]   shiftRegisterNE_26_output_re;
  wire       [23:0]   shiftRegisterNE_26_output_im;
  wire       [23:0]   r2Butterfly_13_out1_re;
  wire       [23:0]   r2Butterfly_13_out1_im;
  wire       [23:0]   r2Butterfly_13_out2_re;
  wire       [23:0]   r2Butterfly_13_out2_im;
  wire       [23:0]   shiftRegisterNE_27_output_re;
  wire       [23:0]   shiftRegisterNE_27_output_im;
  wire       [23:0]   r2Switch_13_out1_re;
  wire       [23:0]   r2Switch_13_out1_im;
  wire       [23:0]   r2Switch_13_out2_re;
  wire       [23:0]   r2Switch_13_out2_im;
  wire       [23:0]   shiftRegisterNE_28_output_re;
  wire       [23:0]   shiftRegisterNE_28_output_im;
  wire       [23:0]   r2Butterfly_14_out1_re;
  wire       [23:0]   r2Butterfly_14_out1_im;
  wire       [23:0]   r2Butterfly_14_out2_re;
  wire       [23:0]   r2Butterfly_14_out2_im;
  wire       [23:0]   shiftRegisterNE_29_output_re;
  wire       [23:0]   shiftRegisterNE_29_output_im;
  wire       [23:0]   r2Switch_14_out1_re;
  wire       [23:0]   r2Switch_14_out1_im;
  wire       [23:0]   r2Switch_14_out2_re;
  wire       [23:0]   r2Switch_14_out2_im;
  wire       [23:0]   shiftRegisterNE_30_output_re;
  wire       [23:0]   shiftRegisterNE_30_output_im;
  wire       [23:0]   r2Butterfly_15_out1_re;
  wire       [23:0]   r2Butterfly_15_out1_im;
  wire       [23:0]   r2Butterfly_15_out2_re;
  wire       [23:0]   r2Butterfly_15_out2_im;
  wire       [23:0]   shiftRegisterNE_31_output_re;
  wire       [23:0]   shiftRegisterNE_31_output_im;
  wire       [23:0]   r2Switch_15_out1_re;
  wire       [23:0]   r2Switch_15_out1_im;
  wire       [23:0]   r2Switch_15_out2_re;
  wire       [23:0]   r2Switch_15_out2_im;
  wire       [23:0]   shiftRegisterNE_32_output_re;
  wire       [23:0]   shiftRegisterNE_32_output_im;
  wire       [23:0]   r2Butterfly_16_out1_re;
  wire       [23:0]   r2Butterfly_16_out1_im;
  wire       [23:0]   r2Butterfly_16_out2_re;
  wire       [23:0]   r2Butterfly_16_out2_im;
  wire       [23:0]   shiftRegisterNE_33_output_re;
  wire       [23:0]   shiftRegisterNE_33_output_im;
  wire       [23:0]   r2Switch_16_out1_re;
  wire       [23:0]   r2Switch_16_out1_im;
  wire       [23:0]   r2Switch_16_out2_re;
  wire       [23:0]   r2Switch_16_out2_im;
  wire       [23:0]   shiftRegisterNE_34_output_re;
  wire       [23:0]   shiftRegisterNE_34_output_im;
  wire       [23:0]   r2Butterfly_17_out1_re;
  wire       [23:0]   r2Butterfly_17_out1_im;
  wire       [23:0]   r2Butterfly_17_out2_re;
  wire       [23:0]   r2Butterfly_17_out2_im;
  wire       [23:0]   shiftRegisterNE_35_output_re;
  wire       [23:0]   shiftRegisterNE_35_output_im;
  wire       [23:0]   r2Switch_17_out1_re;
  wire       [23:0]   r2Switch_17_out1_im;
  wire       [23:0]   r2Switch_17_out2_re;
  wire       [23:0]   r2Switch_17_out2_im;
  wire       [23:0]   shiftRegisterNE_36_output_re;
  wire       [23:0]   shiftRegisterNE_36_output_im;
  wire       [23:0]   r2Butterfly_18_out1_re;
  wire       [23:0]   r2Butterfly_18_out1_im;
  wire       [23:0]   r2Butterfly_18_out2_re;
  wire       [23:0]   r2Butterfly_18_out2_im;
  wire       [23:0]   shiftRegisterNE_37_output_re;
  wire       [23:0]   shiftRegisterNE_37_output_im;
  wire       [23:0]   r2Switch_18_out1_re;
  wire       [23:0]   r2Switch_18_out1_im;
  wire       [23:0]   r2Switch_18_out2_re;
  wire       [23:0]   r2Switch_18_out2_im;
  wire       [23:0]   shiftRegisterNE_38_output_re;
  wire       [23:0]   shiftRegisterNE_38_output_im;
  wire       [23:0]   r2Butterfly_19_out1_re;
  wire       [23:0]   r2Butterfly_19_out1_im;
  wire       [23:0]   r2Butterfly_19_out2_re;
  wire       [23:0]   r2Butterfly_19_out2_im;
  wire       [23:0]   shiftRegisterNE_39_output_re;
  wire       [23:0]   shiftRegisterNE_39_output_im;
  wire       [23:0]   r2Switch_19_out1_re;
  wire       [23:0]   r2Switch_19_out1_im;
  wire       [23:0]   r2Switch_19_out2_re;
  wire       [23:0]   r2Switch_19_out2_im;
  wire                reorder_1_sorted_valid;
  wire                reorder_1_sorted_payload_last;
  wire       [23:0]   reorder_1_sorted_payload_fragment_re;
  wire       [23:0]   reorder_1_sorted_payload_fragment_im;
  wire       [11:0]   _zz_cnt;
  wire                _zz__zz_1_port;
  wire                _zz__zz_wn_re_2;
  wire       [23:0]   _zz__zz_wn_re_1;
  wire       [23:0]   _zz__zz_wn_im;
  wire       [23:0]   _zz_wn_im_10;
  wire       [23:0]   _zz_wn_im_11;
  wire                _zz__zz_2_port;
  wire                _zz__zz_wn_re_5;
  wire       [23:0]   _zz__zz_wn_re_4;
  wire       [23:0]   _zz__zz_wn_im_1;
  wire       [23:0]   _zz_wn_im_12;
  wire       [23:0]   _zz_wn_im_13;
  wire                _zz__zz_3_port;
  wire                _zz__zz_wn_re_8;
  wire       [23:0]   _zz__zz_wn_re_7;
  wire       [23:0]   _zz__zz_wn_im_2;
  wire       [23:0]   _zz_wn_im_14;
  wire       [23:0]   _zz_wn_im_15;
  wire                _zz__zz_4_port;
  wire                _zz__zz_wn_re_11;
  wire       [23:0]   _zz__zz_wn_re_10;
  wire       [23:0]   _zz__zz_wn_im_3;
  wire       [23:0]   _zz_wn_im_16;
  wire       [23:0]   _zz_wn_im_17;
  wire                _zz__zz_5_port;
  wire                _zz__zz_wn_re_14;
  wire       [23:0]   _zz__zz_wn_re_13;
  wire       [23:0]   _zz__zz_wn_im_4;
  wire       [23:0]   _zz_wn_im_18;
  wire       [23:0]   _zz_wn_im_19;
  wire                _zz__zz_6_port;
  wire                _zz__zz_wn_re_17;
  wire       [23:0]   _zz__zz_wn_re_16;
  wire       [23:0]   _zz__zz_wn_im_5;
  wire       [23:0]   _zz_wn_im_20;
  wire       [23:0]   _zz_wn_im_21;
  wire                _zz__zz_7_port;
  wire                _zz__zz_wn_re_20;
  wire       [23:0]   _zz__zz_wn_re_19;
  wire       [23:0]   _zz__zz_wn_im_6;
  wire       [23:0]   _zz_wn_im_22;
  wire       [23:0]   _zz_wn_im_23;
  wire                _zz__zz_8_port;
  wire                _zz__zz_wn_re_23;
  wire       [23:0]   _zz__zz_wn_re_22;
  wire       [23:0]   _zz__zz_wn_im_7;
  wire       [23:0]   _zz_wn_im_24;
  wire       [23:0]   _zz_wn_im_25;
  wire                _zz__zz_9_port;
  wire                _zz__zz_wn_re_26;
  wire       [23:0]   _zz__zz_wn_re_25;
  wire       [23:0]   _zz__zz_wn_im_8;
  wire       [23:0]   _zz_wn_im_26;
  wire       [23:0]   _zz_wn_im_27;
  wire                _zz__zz_10_port;
  wire                _zz__zz_wn_re_29;
  wire       [23:0]   _zz__zz_wn_re_28;
  wire       [23:0]   _zz__zz_wn_im_9;
  wire       [23:0]   _zz_wn_im_28;
  wire       [23:0]   _zz_wn_im_29;
  wire       [23:0]   _zz_result_out1_re;
  wire       [12:0]   _zz_result_out1_re_1;
  wire       [23:0]   _zz_result_out1_im;
  wire       [12:0]   _zz_result_out1_im_1;
  wire       [23:0]   _zz_result_out2_re;
  wire       [12:0]   _zz_result_out2_re_1;
  wire       [23:0]   _zz_result_out2_im;
  wire       [12:0]   _zz_result_out2_im_1;
  reg        [11:0]   cnt;
  wire                raw_data_fire;
  wire                when_R2MDC_l20;
  wire       [23:0]   out0_buf_0_re;
  wire       [23:0]   out0_buf_0_im;
  wire       [23:0]   out0_buf_1_re;
  wire       [23:0]   out0_buf_1_im;
  wire       [23:0]   out0_buf_2_re;
  wire       [23:0]   out0_buf_2_im;
  wire       [23:0]   out0_buf_3_re;
  wire       [23:0]   out0_buf_3_im;
  wire       [23:0]   out0_buf_4_re;
  wire       [23:0]   out0_buf_4_im;
  wire       [23:0]   out0_buf_5_re;
  wire       [23:0]   out0_buf_5_im;
  wire       [23:0]   out0_buf_6_re;
  wire       [23:0]   out0_buf_6_im;
  wire       [23:0]   out0_buf_7_re;
  wire       [23:0]   out0_buf_7_im;
  wire       [23:0]   out0_buf_8_re;
  wire       [23:0]   out0_buf_8_im;
  wire       [23:0]   out0_buf_9_re;
  wire       [23:0]   out0_buf_9_im;
  wire       [23:0]   out0_buf_10_re;
  wire       [23:0]   out0_buf_10_im;
  wire       [23:0]   out0_buf_11_re;
  wire       [23:0]   out0_buf_11_im;
  wire       [23:0]   out1_buf_0_re;
  wire       [23:0]   out1_buf_0_im;
  wire       [23:0]   out1_buf_1_re;
  wire       [23:0]   out1_buf_1_im;
  wire       [23:0]   out1_buf_2_re;
  wire       [23:0]   out1_buf_2_im;
  wire       [23:0]   out1_buf_3_re;
  wire       [23:0]   out1_buf_3_im;
  wire       [23:0]   out1_buf_4_re;
  wire       [23:0]   out1_buf_4_im;
  wire       [23:0]   out1_buf_5_re;
  wire       [23:0]   out1_buf_5_im;
  wire       [23:0]   out1_buf_6_re;
  wire       [23:0]   out1_buf_6_im;
  wire       [23:0]   out1_buf_7_re;
  wire       [23:0]   out1_buf_7_im;
  wire       [23:0]   out1_buf_8_re;
  wire       [23:0]   out1_buf_8_im;
  wire       [23:0]   out1_buf_9_re;
  wire       [23:0]   out1_buf_9_im;
  wire       [23:0]   out1_buf_10_re;
  wire       [23:0]   out1_buf_10_im;
  wire       [23:0]   out1_buf_11_re;
  wire       [23:0]   out1_buf_11_im;
  wire       [11:0]   cnt_p1;
  wire       [9:0]    _zz_wn_re;
  wire       [23:0]   _zz_wn_re_1;
  wire       [23:0]   _zz_wn_im;
  wire       [47:0]   _zz_wn_re_2;
  wire       [8:0]    _zz_wn_re_3;
  wire       [23:0]   _zz_wn_re_4;
  wire       [23:0]   _zz_wn_im_1;
  wire       [47:0]   _zz_wn_re_5;
  wire       [7:0]    _zz_wn_re_6;
  wire       [23:0]   _zz_wn_re_7;
  wire       [23:0]   _zz_wn_im_2;
  wire       [47:0]   _zz_wn_re_8;
  wire       [6:0]    _zz_wn_re_9;
  wire       [23:0]   _zz_wn_re_10;
  wire       [23:0]   _zz_wn_im_3;
  wire       [47:0]   _zz_wn_re_11;
  wire       [5:0]    _zz_wn_re_12;
  wire       [23:0]   _zz_wn_re_13;
  wire       [23:0]   _zz_wn_im_4;
  wire       [47:0]   _zz_wn_re_14;
  wire       [4:0]    _zz_wn_re_15;
  wire       [23:0]   _zz_wn_re_16;
  wire       [23:0]   _zz_wn_im_5;
  wire       [47:0]   _zz_wn_re_17;
  wire       [3:0]    _zz_wn_re_18;
  wire       [23:0]   _zz_wn_re_19;
  wire       [23:0]   _zz_wn_im_6;
  wire       [47:0]   _zz_wn_re_20;
  wire       [2:0]    _zz_wn_re_21;
  wire       [23:0]   _zz_wn_re_22;
  wire       [23:0]   _zz_wn_im_7;
  wire       [47:0]   _zz_wn_re_23;
  wire       [1:0]    _zz_wn_re_24;
  wire       [23:0]   _zz_wn_re_25;
  wire       [23:0]   _zz_wn_im_8;
  wire       [47:0]   _zz_wn_re_26;
  wire       [0:0]    _zz_wn_re_27;
  wire       [23:0]   _zz_wn_re_28;
  wire       [23:0]   _zz_wn_im_9;
  wire       [47:0]   _zz_wn_re_29;
  reg        [23:0]   out1D1_re;
  reg        [23:0]   out1D1_im;
  wire       [23:0]   result_out1_re;
  wire       [23:0]   result_out1_im;
  wire       [23:0]   result_out2_re;
  wire       [23:0]   result_out2_im;
  reg        [23:0]   result_out1_regNext_re;
  reg        [23:0]   result_out1_regNext_im;
  reg        [23:0]   result_out2_regNext_re;
  reg        [23:0]   result_out2_regNext_im;
  (* rom_style = "block" *) reg [47:0] _zz_1 [0:1023];
  (* rom_style = "block" *) reg [47:0] _zz_2 [0:511];
  (* rom_style = "block" *) reg [47:0] _zz_3 [0:255];
  (* rom_style = "block" *) reg [47:0] _zz_4 [0:127];
  (* rom_style = "block" *) reg [47:0] _zz_5 [0:63];
  (* rom_style = "block" *) reg [47:0] _zz_6 [0:31];
  (* rom_style = "block" *) reg [47:0] _zz_7 [0:15];
  (* rom_style = "block" *) reg [47:0] _zz_8 [0:7];
  (* rom_style = "block" *) reg [47:0] _zz_9 [0:3];
  (* rom_style = "block" *) reg [47:0] _zz_10 [0:1];

  assign _zz_cnt = (cnt + 12'h001);
  assign _zz__zz_wn_re_1 = _zz_wn_re_2[23 : 0];
  assign _zz__zz_wn_im = _zz_wn_re_2[47 : 24];
  assign _zz_wn_im_10 = ($signed(_zz_wn_im_11) - $signed(_zz_wn_im));
  assign _zz_wn_im_11 = 24'h0;
  assign _zz__zz_wn_re_4 = _zz_wn_re_5[23 : 0];
  assign _zz__zz_wn_im_1 = _zz_wn_re_5[47 : 24];
  assign _zz_wn_im_12 = ($signed(_zz_wn_im_13) - $signed(_zz_wn_im_1));
  assign _zz_wn_im_13 = 24'h0;
  assign _zz__zz_wn_re_7 = _zz_wn_re_8[23 : 0];
  assign _zz__zz_wn_im_2 = _zz_wn_re_8[47 : 24];
  assign _zz_wn_im_14 = ($signed(_zz_wn_im_15) - $signed(_zz_wn_im_2));
  assign _zz_wn_im_15 = 24'h0;
  assign _zz__zz_wn_re_10 = _zz_wn_re_11[23 : 0];
  assign _zz__zz_wn_im_3 = _zz_wn_re_11[47 : 24];
  assign _zz_wn_im_16 = ($signed(_zz_wn_im_17) - $signed(_zz_wn_im_3));
  assign _zz_wn_im_17 = 24'h0;
  assign _zz__zz_wn_re_13 = _zz_wn_re_14[23 : 0];
  assign _zz__zz_wn_im_4 = _zz_wn_re_14[47 : 24];
  assign _zz_wn_im_18 = ($signed(_zz_wn_im_19) - $signed(_zz_wn_im_4));
  assign _zz_wn_im_19 = 24'h0;
  assign _zz__zz_wn_re_16 = _zz_wn_re_17[23 : 0];
  assign _zz__zz_wn_im_5 = _zz_wn_re_17[47 : 24];
  assign _zz_wn_im_20 = ($signed(_zz_wn_im_21) - $signed(_zz_wn_im_5));
  assign _zz_wn_im_21 = 24'h0;
  assign _zz__zz_wn_re_19 = _zz_wn_re_20[23 : 0];
  assign _zz__zz_wn_im_6 = _zz_wn_re_20[47 : 24];
  assign _zz_wn_im_22 = ($signed(_zz_wn_im_23) - $signed(_zz_wn_im_6));
  assign _zz_wn_im_23 = 24'h0;
  assign _zz__zz_wn_re_22 = _zz_wn_re_23[23 : 0];
  assign _zz__zz_wn_im_7 = _zz_wn_re_23[47 : 24];
  assign _zz_wn_im_24 = ($signed(_zz_wn_im_25) - $signed(_zz_wn_im_7));
  assign _zz_wn_im_25 = 24'h0;
  assign _zz__zz_wn_re_25 = _zz_wn_re_26[23 : 0];
  assign _zz__zz_wn_im_8 = _zz_wn_re_26[47 : 24];
  assign _zz_wn_im_26 = ($signed(_zz_wn_im_27) - $signed(_zz_wn_im_8));
  assign _zz_wn_im_27 = 24'h0;
  assign _zz__zz_wn_re_28 = _zz_wn_re_29[23 : 0];
  assign _zz__zz_wn_im_9 = _zz_wn_re_29[47 : 24];
  assign _zz_wn_im_28 = ($signed(_zz_wn_im_29) - $signed(_zz_wn_im_9));
  assign _zz_wn_im_29 = 24'h0;
  assign _zz_result_out1_re_1 = (out0_buf_11_re >>> 11);
  assign _zz_result_out1_re = {{11{_zz_result_out1_re_1[12]}}, _zz_result_out1_re_1};
  assign _zz_result_out1_im_1 = (out0_buf_11_im >>> 11);
  assign _zz_result_out1_im = {{11{_zz_result_out1_im_1[12]}}, _zz_result_out1_im_1};
  assign _zz_result_out2_re_1 = (out1_buf_11_re >>> 11);
  assign _zz_result_out2_re = {{11{_zz_result_out2_re_1[12]}}, _zz_result_out2_re_1};
  assign _zz_result_out2_im_1 = (out1_buf_11_im >>> 11);
  assign _zz_result_out2_im = {{11{_zz_result_out2_im_1[12]}}, _zz_result_out2_im_1};
  assign _zz__zz_wn_re_2 = 1'b1;
  assign _zz__zz_wn_re_5 = 1'b1;
  assign _zz__zz_wn_re_8 = 1'b1;
  assign _zz__zz_wn_re_11 = 1'b1;
  assign _zz__zz_wn_re_14 = 1'b1;
  assign _zz__zz_wn_re_17 = 1'b1;
  assign _zz__zz_wn_re_20 = 1'b1;
  assign _zz__zz_wn_re_23 = 1'b1;
  assign _zz__zz_wn_re_26 = 1'b1;
  assign _zz__zz_wn_re_29 = 1'b1;
  initial begin
    $readmemb("R2MDC.v_toplevel__zz_1.bin",_zz_1);
  end
  always @(posedge clk) begin
    if(_zz__zz_wn_re_2) begin
      _zz__zz_1_port0 <= _zz_1[_zz_wn_re];
    end
  end

  initial begin
    $readmemb("R2MDC.v_toplevel__zz_2.bin",_zz_2);
  end
  always @(posedge clk) begin
    if(_zz__zz_wn_re_5) begin
      _zz__zz_2_port0 <= _zz_2[_zz_wn_re_3];
    end
  end

  initial begin
    $readmemb("R2MDC.v_toplevel__zz_3.bin",_zz_3);
  end
  always @(posedge clk) begin
    if(_zz__zz_wn_re_8) begin
      _zz__zz_3_port0 <= _zz_3[_zz_wn_re_6];
    end
  end

  initial begin
    $readmemb("R2MDC.v_toplevel__zz_4.bin",_zz_4);
  end
  always @(posedge clk) begin
    if(_zz__zz_wn_re_11) begin
      _zz__zz_4_port0 <= _zz_4[_zz_wn_re_9];
    end
  end

  initial begin
    $readmemb("R2MDC.v_toplevel__zz_5.bin",_zz_5);
  end
  always @(posedge clk) begin
    if(_zz__zz_wn_re_14) begin
      _zz__zz_5_port0 <= _zz_5[_zz_wn_re_12];
    end
  end

  initial begin
    $readmemb("R2MDC.v_toplevel__zz_6.bin",_zz_6);
  end
  always @(posedge clk) begin
    if(_zz__zz_wn_re_17) begin
      _zz__zz_6_port0 <= _zz_6[_zz_wn_re_15];
    end
  end

  initial begin
    $readmemb("R2MDC.v_toplevel__zz_7.bin",_zz_7);
  end
  always @(posedge clk) begin
    if(_zz__zz_wn_re_20) begin
      _zz__zz_7_port0 <= _zz_7[_zz_wn_re_18];
    end
  end

  initial begin
    $readmemb("R2MDC.v_toplevel__zz_8.bin",_zz_8);
  end
  always @(posedge clk) begin
    if(_zz__zz_wn_re_23) begin
      _zz__zz_8_port0 <= _zz_8[_zz_wn_re_21];
    end
  end

  initial begin
    $readmemb("R2MDC.v_toplevel__zz_9.bin",_zz_9);
  end
  always @(posedge clk) begin
    if(_zz__zz_wn_re_26) begin
      _zz__zz_9_port0 <= _zz_9[_zz_wn_re_24];
    end
  end

  initial begin
    $readmemb("R2MDC.v_toplevel__zz_10.bin",_zz_10);
  end
  always @(posedge clk) begin
    if(_zz__zz_wn_re_29) begin
      _zz__zz_10_port0 <= _zz_10[_zz_wn_re_27];
    end
  end

  ShiftRegisterNE shiftRegisterNE_20 (
    .input_re     (out0_buf_0_re                 ), //i
    .input_im     (out0_buf_0_im                 ), //i
    .output_re    (shiftRegisterNE_20_output_re  ), //o
    .output_im    (shiftRegisterNE_20_output_im  ), //o
    .clk          (clk                           ), //i
    .reset        (reset                         )  //i
  );
  R2Butterfly r2Butterfly_10 (
    .in1_re     (shiftRegisterNE_20_output_re  ), //i
    .in1_im     (shiftRegisterNE_20_output_im  ), //i
    .in2_re     (out1_buf_0_re                 ), //i
    .in2_im     (out1_buf_0_im                 ), //i
    .wn_re      (r2Butterfly_10_wn_re          ), //i
    .wn_im      (r2Butterfly_10_wn_im          ), //i
    .out1_re    (r2Butterfly_10_out1_re        ), //o
    .out1_im    (r2Butterfly_10_out1_im        ), //o
    .out2_re    (r2Butterfly_10_out2_re        ), //o
    .out2_im    (r2Butterfly_10_out2_im        )  //o
  );
  ShiftRegisterNE_1 shiftRegisterNE_21 (
    .input_re     (r2Butterfly_10_out2_re        ), //i
    .input_im     (r2Butterfly_10_out2_im        ), //i
    .output_re    (shiftRegisterNE_21_output_re  ), //o
    .output_im    (shiftRegisterNE_21_output_im  ), //o
    .clk          (clk                           ), //i
    .reset        (reset                         )  //i
  );
  R2Switch r2Switch_10 (
    .in1_re     (r2Butterfly_10_out1_re        ), //i
    .in1_im     (r2Butterfly_10_out1_im        ), //i
    .in2_re     (shiftRegisterNE_21_output_re  ), //i
    .in2_im     (shiftRegisterNE_21_output_im  ), //i
    .sel        (r2Switch_10_sel               ), //i
    .out1_re    (r2Switch_10_out1_re           ), //o
    .out1_im    (r2Switch_10_out1_im           ), //o
    .out2_re    (r2Switch_10_out2_re           ), //o
    .out2_im    (r2Switch_10_out2_im           )  //o
  );
  ShiftRegisterNE_1 shiftRegisterNE_22 (
    .input_re     (out0_buf_1_re                 ), //i
    .input_im     (out0_buf_1_im                 ), //i
    .output_re    (shiftRegisterNE_22_output_re  ), //o
    .output_im    (shiftRegisterNE_22_output_im  ), //o
    .clk          (clk                           ), //i
    .reset        (reset                         )  //i
  );
  R2Butterfly r2Butterfly_11 (
    .in1_re     (shiftRegisterNE_22_output_re  ), //i
    .in1_im     (shiftRegisterNE_22_output_im  ), //i
    .in2_re     (out1_buf_1_re                 ), //i
    .in2_im     (out1_buf_1_im                 ), //i
    .wn_re      (r2Butterfly_11_wn_re          ), //i
    .wn_im      (r2Butterfly_11_wn_im          ), //i
    .out1_re    (r2Butterfly_11_out1_re        ), //o
    .out1_im    (r2Butterfly_11_out1_im        ), //o
    .out2_re    (r2Butterfly_11_out2_re        ), //o
    .out2_im    (r2Butterfly_11_out2_im        )  //o
  );
  ShiftRegisterNE_3 shiftRegisterNE_23 (
    .input_re     (r2Butterfly_11_out2_re        ), //i
    .input_im     (r2Butterfly_11_out2_im        ), //i
    .output_re    (shiftRegisterNE_23_output_re  ), //o
    .output_im    (shiftRegisterNE_23_output_im  ), //o
    .clk          (clk                           ), //i
    .reset        (reset                         )  //i
  );
  R2Switch r2Switch_11 (
    .in1_re     (r2Butterfly_11_out1_re        ), //i
    .in1_im     (r2Butterfly_11_out1_im        ), //i
    .in2_re     (shiftRegisterNE_23_output_re  ), //i
    .in2_im     (shiftRegisterNE_23_output_im  ), //i
    .sel        (r2Switch_11_sel               ), //i
    .out1_re    (r2Switch_11_out1_re           ), //o
    .out1_im    (r2Switch_11_out1_im           ), //o
    .out2_re    (r2Switch_11_out2_re           ), //o
    .out2_im    (r2Switch_11_out2_im           )  //o
  );
  ShiftRegisterNE_3 shiftRegisterNE_24 (
    .input_re     (out0_buf_2_re                 ), //i
    .input_im     (out0_buf_2_im                 ), //i
    .output_re    (shiftRegisterNE_24_output_re  ), //o
    .output_im    (shiftRegisterNE_24_output_im  ), //o
    .clk          (clk                           ), //i
    .reset        (reset                         )  //i
  );
  R2Butterfly r2Butterfly_12 (
    .in1_re     (shiftRegisterNE_24_output_re  ), //i
    .in1_im     (shiftRegisterNE_24_output_im  ), //i
    .in2_re     (out1_buf_2_re                 ), //i
    .in2_im     (out1_buf_2_im                 ), //i
    .wn_re      (r2Butterfly_12_wn_re          ), //i
    .wn_im      (r2Butterfly_12_wn_im          ), //i
    .out1_re    (r2Butterfly_12_out1_re        ), //o
    .out1_im    (r2Butterfly_12_out1_im        ), //o
    .out2_re    (r2Butterfly_12_out2_re        ), //o
    .out2_im    (r2Butterfly_12_out2_im        )  //o
  );
  ShiftRegisterNE_5 shiftRegisterNE_25 (
    .input_re     (r2Butterfly_12_out2_re        ), //i
    .input_im     (r2Butterfly_12_out2_im        ), //i
    .output_re    (shiftRegisterNE_25_output_re  ), //o
    .output_im    (shiftRegisterNE_25_output_im  ), //o
    .clk          (clk                           ), //i
    .reset        (reset                         )  //i
  );
  R2Switch r2Switch_12 (
    .in1_re     (r2Butterfly_12_out1_re        ), //i
    .in1_im     (r2Butterfly_12_out1_im        ), //i
    .in2_re     (shiftRegisterNE_25_output_re  ), //i
    .in2_im     (shiftRegisterNE_25_output_im  ), //i
    .sel        (r2Switch_12_sel               ), //i
    .out1_re    (r2Switch_12_out1_re           ), //o
    .out1_im    (r2Switch_12_out1_im           ), //o
    .out2_re    (r2Switch_12_out2_re           ), //o
    .out2_im    (r2Switch_12_out2_im           )  //o
  );
  ShiftRegisterNE_5 shiftRegisterNE_26 (
    .input_re     (out0_buf_3_re                 ), //i
    .input_im     (out0_buf_3_im                 ), //i
    .output_re    (shiftRegisterNE_26_output_re  ), //o
    .output_im    (shiftRegisterNE_26_output_im  ), //o
    .clk          (clk                           ), //i
    .reset        (reset                         )  //i
  );
  R2Butterfly r2Butterfly_13 (
    .in1_re     (shiftRegisterNE_26_output_re  ), //i
    .in1_im     (shiftRegisterNE_26_output_im  ), //i
    .in2_re     (out1_buf_3_re                 ), //i
    .in2_im     (out1_buf_3_im                 ), //i
    .wn_re      (r2Butterfly_13_wn_re          ), //i
    .wn_im      (r2Butterfly_13_wn_im          ), //i
    .out1_re    (r2Butterfly_13_out1_re        ), //o
    .out1_im    (r2Butterfly_13_out1_im        ), //o
    .out2_re    (r2Butterfly_13_out2_re        ), //o
    .out2_im    (r2Butterfly_13_out2_im        )  //o
  );
  ShiftRegisterNE_7 shiftRegisterNE_27 (
    .input_re     (r2Butterfly_13_out2_re        ), //i
    .input_im     (r2Butterfly_13_out2_im        ), //i
    .output_re    (shiftRegisterNE_27_output_re  ), //o
    .output_im    (shiftRegisterNE_27_output_im  ), //o
    .clk          (clk                           ), //i
    .reset        (reset                         )  //i
  );
  R2Switch r2Switch_13 (
    .in1_re     (r2Butterfly_13_out1_re        ), //i
    .in1_im     (r2Butterfly_13_out1_im        ), //i
    .in2_re     (shiftRegisterNE_27_output_re  ), //i
    .in2_im     (shiftRegisterNE_27_output_im  ), //i
    .sel        (r2Switch_13_sel               ), //i
    .out1_re    (r2Switch_13_out1_re           ), //o
    .out1_im    (r2Switch_13_out1_im           ), //o
    .out2_re    (r2Switch_13_out2_re           ), //o
    .out2_im    (r2Switch_13_out2_im           )  //o
  );
  ShiftRegisterNE_7 shiftRegisterNE_28 (
    .input_re     (out0_buf_4_re                 ), //i
    .input_im     (out0_buf_4_im                 ), //i
    .output_re    (shiftRegisterNE_28_output_re  ), //o
    .output_im    (shiftRegisterNE_28_output_im  ), //o
    .clk          (clk                           ), //i
    .reset        (reset                         )  //i
  );
  R2Butterfly r2Butterfly_14 (
    .in1_re     (shiftRegisterNE_28_output_re  ), //i
    .in1_im     (shiftRegisterNE_28_output_im  ), //i
    .in2_re     (out1_buf_4_re                 ), //i
    .in2_im     (out1_buf_4_im                 ), //i
    .wn_re      (r2Butterfly_14_wn_re          ), //i
    .wn_im      (r2Butterfly_14_wn_im          ), //i
    .out1_re    (r2Butterfly_14_out1_re        ), //o
    .out1_im    (r2Butterfly_14_out1_im        ), //o
    .out2_re    (r2Butterfly_14_out2_re        ), //o
    .out2_im    (r2Butterfly_14_out2_im        )  //o
  );
  ShiftRegisterNE_9 shiftRegisterNE_29 (
    .input_re     (r2Butterfly_14_out2_re        ), //i
    .input_im     (r2Butterfly_14_out2_im        ), //i
    .output_re    (shiftRegisterNE_29_output_re  ), //o
    .output_im    (shiftRegisterNE_29_output_im  ), //o
    .clk          (clk                           ), //i
    .reset        (reset                         )  //i
  );
  R2Switch r2Switch_14 (
    .in1_re     (r2Butterfly_14_out1_re        ), //i
    .in1_im     (r2Butterfly_14_out1_im        ), //i
    .in2_re     (shiftRegisterNE_29_output_re  ), //i
    .in2_im     (shiftRegisterNE_29_output_im  ), //i
    .sel        (r2Switch_14_sel               ), //i
    .out1_re    (r2Switch_14_out1_re           ), //o
    .out1_im    (r2Switch_14_out1_im           ), //o
    .out2_re    (r2Switch_14_out2_re           ), //o
    .out2_im    (r2Switch_14_out2_im           )  //o
  );
  ShiftRegisterNE_9 shiftRegisterNE_30 (
    .input_re     (out0_buf_5_re                 ), //i
    .input_im     (out0_buf_5_im                 ), //i
    .output_re    (shiftRegisterNE_30_output_re  ), //o
    .output_im    (shiftRegisterNE_30_output_im  ), //o
    .clk          (clk                           ), //i
    .reset        (reset                         )  //i
  );
  R2Butterfly r2Butterfly_15 (
    .in1_re     (shiftRegisterNE_30_output_re  ), //i
    .in1_im     (shiftRegisterNE_30_output_im  ), //i
    .in2_re     (out1_buf_5_re                 ), //i
    .in2_im     (out1_buf_5_im                 ), //i
    .wn_re      (r2Butterfly_15_wn_re          ), //i
    .wn_im      (r2Butterfly_15_wn_im          ), //i
    .out1_re    (r2Butterfly_15_out1_re        ), //o
    .out1_im    (r2Butterfly_15_out1_im        ), //o
    .out2_re    (r2Butterfly_15_out2_re        ), //o
    .out2_im    (r2Butterfly_15_out2_im        )  //o
  );
  ShiftRegisterNE_11 shiftRegisterNE_31 (
    .input_re     (r2Butterfly_15_out2_re        ), //i
    .input_im     (r2Butterfly_15_out2_im        ), //i
    .output_re    (shiftRegisterNE_31_output_re  ), //o
    .output_im    (shiftRegisterNE_31_output_im  ), //o
    .clk          (clk                           ), //i
    .reset        (reset                         )  //i
  );
  R2Switch r2Switch_15 (
    .in1_re     (r2Butterfly_15_out1_re        ), //i
    .in1_im     (r2Butterfly_15_out1_im        ), //i
    .in2_re     (shiftRegisterNE_31_output_re  ), //i
    .in2_im     (shiftRegisterNE_31_output_im  ), //i
    .sel        (r2Switch_15_sel               ), //i
    .out1_re    (r2Switch_15_out1_re           ), //o
    .out1_im    (r2Switch_15_out1_im           ), //o
    .out2_re    (r2Switch_15_out2_re           ), //o
    .out2_im    (r2Switch_15_out2_im           )  //o
  );
  ShiftRegisterNE_11 shiftRegisterNE_32 (
    .input_re     (out0_buf_6_re                 ), //i
    .input_im     (out0_buf_6_im                 ), //i
    .output_re    (shiftRegisterNE_32_output_re  ), //o
    .output_im    (shiftRegisterNE_32_output_im  ), //o
    .clk          (clk                           ), //i
    .reset        (reset                         )  //i
  );
  R2Butterfly r2Butterfly_16 (
    .in1_re     (shiftRegisterNE_32_output_re  ), //i
    .in1_im     (shiftRegisterNE_32_output_im  ), //i
    .in2_re     (out1_buf_6_re                 ), //i
    .in2_im     (out1_buf_6_im                 ), //i
    .wn_re      (r2Butterfly_16_wn_re          ), //i
    .wn_im      (r2Butterfly_16_wn_im          ), //i
    .out1_re    (r2Butterfly_16_out1_re        ), //o
    .out1_im    (r2Butterfly_16_out1_im        ), //o
    .out2_re    (r2Butterfly_16_out2_re        ), //o
    .out2_im    (r2Butterfly_16_out2_im        )  //o
  );
  ShiftRegisterNE_13 shiftRegisterNE_33 (
    .input_re     (r2Butterfly_16_out2_re        ), //i
    .input_im     (r2Butterfly_16_out2_im        ), //i
    .output_re    (shiftRegisterNE_33_output_re  ), //o
    .output_im    (shiftRegisterNE_33_output_im  ), //o
    .clk          (clk                           ), //i
    .reset        (reset                         )  //i
  );
  R2Switch r2Switch_16 (
    .in1_re     (r2Butterfly_16_out1_re        ), //i
    .in1_im     (r2Butterfly_16_out1_im        ), //i
    .in2_re     (shiftRegisterNE_33_output_re  ), //i
    .in2_im     (shiftRegisterNE_33_output_im  ), //i
    .sel        (r2Switch_16_sel               ), //i
    .out1_re    (r2Switch_16_out1_re           ), //o
    .out1_im    (r2Switch_16_out1_im           ), //o
    .out2_re    (r2Switch_16_out2_re           ), //o
    .out2_im    (r2Switch_16_out2_im           )  //o
  );
  ShiftRegisterNE_13 shiftRegisterNE_34 (
    .input_re     (out0_buf_7_re                 ), //i
    .input_im     (out0_buf_7_im                 ), //i
    .output_re    (shiftRegisterNE_34_output_re  ), //o
    .output_im    (shiftRegisterNE_34_output_im  ), //o
    .clk          (clk                           ), //i
    .reset        (reset                         )  //i
  );
  R2Butterfly r2Butterfly_17 (
    .in1_re     (shiftRegisterNE_34_output_re  ), //i
    .in1_im     (shiftRegisterNE_34_output_im  ), //i
    .in2_re     (out1_buf_7_re                 ), //i
    .in2_im     (out1_buf_7_im                 ), //i
    .wn_re      (r2Butterfly_17_wn_re          ), //i
    .wn_im      (r2Butterfly_17_wn_im          ), //i
    .out1_re    (r2Butterfly_17_out1_re        ), //o
    .out1_im    (r2Butterfly_17_out1_im        ), //o
    .out2_re    (r2Butterfly_17_out2_re        ), //o
    .out2_im    (r2Butterfly_17_out2_im        )  //o
  );
  ShiftRegisterNE_15 shiftRegisterNE_35 (
    .input_re     (r2Butterfly_17_out2_re        ), //i
    .input_im     (r2Butterfly_17_out2_im        ), //i
    .output_re    (shiftRegisterNE_35_output_re  ), //o
    .output_im    (shiftRegisterNE_35_output_im  ), //o
    .clk          (clk                           ), //i
    .reset        (reset                         )  //i
  );
  R2Switch r2Switch_17 (
    .in1_re     (r2Butterfly_17_out1_re        ), //i
    .in1_im     (r2Butterfly_17_out1_im        ), //i
    .in2_re     (shiftRegisterNE_35_output_re  ), //i
    .in2_im     (shiftRegisterNE_35_output_im  ), //i
    .sel        (r2Switch_17_sel               ), //i
    .out1_re    (r2Switch_17_out1_re           ), //o
    .out1_im    (r2Switch_17_out1_im           ), //o
    .out2_re    (r2Switch_17_out2_re           ), //o
    .out2_im    (r2Switch_17_out2_im           )  //o
  );
  ShiftRegisterNE_15 shiftRegisterNE_36 (
    .input_re     (out0_buf_8_re                 ), //i
    .input_im     (out0_buf_8_im                 ), //i
    .output_re    (shiftRegisterNE_36_output_re  ), //o
    .output_im    (shiftRegisterNE_36_output_im  ), //o
    .clk          (clk                           ), //i
    .reset        (reset                         )  //i
  );
  R2Butterfly r2Butterfly_18 (
    .in1_re     (shiftRegisterNE_36_output_re  ), //i
    .in1_im     (shiftRegisterNE_36_output_im  ), //i
    .in2_re     (out1_buf_8_re                 ), //i
    .in2_im     (out1_buf_8_im                 ), //i
    .wn_re      (r2Butterfly_18_wn_re          ), //i
    .wn_im      (r2Butterfly_18_wn_im          ), //i
    .out1_re    (r2Butterfly_18_out1_re        ), //o
    .out1_im    (r2Butterfly_18_out1_im        ), //o
    .out2_re    (r2Butterfly_18_out2_re        ), //o
    .out2_im    (r2Butterfly_18_out2_im        )  //o
  );
  ShiftRegisterNE_17 shiftRegisterNE_37 (
    .input_re     (r2Butterfly_18_out2_re        ), //i
    .input_im     (r2Butterfly_18_out2_im        ), //i
    .output_re    (shiftRegisterNE_37_output_re  ), //o
    .output_im    (shiftRegisterNE_37_output_im  ), //o
    .clk          (clk                           ), //i
    .reset        (reset                         )  //i
  );
  R2Switch r2Switch_18 (
    .in1_re     (r2Butterfly_18_out1_re        ), //i
    .in1_im     (r2Butterfly_18_out1_im        ), //i
    .in2_re     (shiftRegisterNE_37_output_re  ), //i
    .in2_im     (shiftRegisterNE_37_output_im  ), //i
    .sel        (r2Switch_18_sel               ), //i
    .out1_re    (r2Switch_18_out1_re           ), //o
    .out1_im    (r2Switch_18_out1_im           ), //o
    .out2_re    (r2Switch_18_out2_re           ), //o
    .out2_im    (r2Switch_18_out2_im           )  //o
  );
  ShiftRegisterNE_17 shiftRegisterNE_38 (
    .input_re     (out0_buf_9_re                 ), //i
    .input_im     (out0_buf_9_im                 ), //i
    .output_re    (shiftRegisterNE_38_output_re  ), //o
    .output_im    (shiftRegisterNE_38_output_im  ), //o
    .clk          (clk                           ), //i
    .reset        (reset                         )  //i
  );
  R2Butterfly r2Butterfly_19 (
    .in1_re     (shiftRegisterNE_38_output_re  ), //i
    .in1_im     (shiftRegisterNE_38_output_im  ), //i
    .in2_re     (out1_buf_9_re                 ), //i
    .in2_im     (out1_buf_9_im                 ), //i
    .wn_re      (r2Butterfly_19_wn_re          ), //i
    .wn_im      (r2Butterfly_19_wn_im          ), //i
    .out1_re    (r2Butterfly_19_out1_re        ), //o
    .out1_im    (r2Butterfly_19_out1_im        ), //o
    .out2_re    (r2Butterfly_19_out2_re        ), //o
    .out2_im    (r2Butterfly_19_out2_im        )  //o
  );
  ShiftRegisterNE_19 shiftRegisterNE_39 (
    .input_re     (r2Butterfly_19_out2_re        ), //i
    .input_im     (r2Butterfly_19_out2_im        ), //i
    .output_re    (shiftRegisterNE_39_output_re  ), //o
    .output_im    (shiftRegisterNE_39_output_im  ), //o
    .clk          (clk                           ), //i
    .reset        (reset                         )  //i
  );
  R2Switch r2Switch_19 (
    .in1_re     (r2Butterfly_19_out1_re        ), //i
    .in1_im     (r2Butterfly_19_out1_im        ), //i
    .in2_re     (shiftRegisterNE_39_output_re  ), //i
    .in2_im     (shiftRegisterNE_39_output_im  ), //i
    .sel        (r2Switch_19_sel               ), //i
    .out1_re    (r2Switch_19_out1_re           ), //o
    .out1_im    (r2Switch_19_out1_im           ), //o
    .out2_re    (r2Switch_19_out2_re           ), //o
    .out2_im    (r2Switch_19_out2_im           )  //o
  );
  Reorder reorder_1 (
    .unsorted_valid                (reorder_1_unsorted_valid              ), //i
    .unsorted_payload_in0_re       (result_out1_regNext_re                ), //i
    .unsorted_payload_in0_im       (result_out1_regNext_im                ), //i
    .unsorted_payload_in1_re       (result_out2_regNext_re                ), //i
    .unsorted_payload_in1_im       (result_out2_regNext_im                ), //i
    .sorted_valid                  (reorder_1_sorted_valid                ), //o
    .sorted_payload_last           (reorder_1_sorted_payload_last         ), //o
    .sorted_payload_fragment_re    (reorder_1_sorted_payload_fragment_re  ), //o
    .sorted_payload_fragment_im    (reorder_1_sorted_payload_fragment_im  ), //o
    .clk                           (clk                                   ), //i
    .reset                         (reset                                 )  //i
  );
  assign raw_data_fire = (raw_data_valid && raw_data_ready);
  assign when_R2MDC_l20 = (raw_data_fire || (12'h800 <= cnt));
  assign raw_data_ready = (cnt < 12'h800);
  assign out0_buf_0_re = raw_data_payload_re;
  assign out0_buf_0_im = raw_data_payload_im;
  assign out1_buf_0_re = raw_data_payload_re;
  assign out1_buf_0_im = raw_data_payload_im;
  assign cnt_p1 = (cnt + 12'h001);
  assign _zz_wn_re = cnt_p1[9 : 0];
  assign _zz_wn_re_2 = _zz__zz_1_port0;
  assign _zz_wn_re_1 = _zz__zz_wn_re_1[23 : 0];
  assign _zz_wn_im = _zz__zz_wn_im[23 : 0];
  assign r2Butterfly_10_wn_re = (mode ? _zz_wn_re_1 : _zz_wn_re_1);
  assign r2Butterfly_10_wn_im = (mode ? _zz_wn_im : _zz_wn_im_10);
  assign r2Switch_10_sel = cnt[9];
  assign out0_buf_1_re = r2Switch_10_out1_re;
  assign out0_buf_1_im = r2Switch_10_out1_im;
  assign out1_buf_1_re = r2Switch_10_out2_re;
  assign out1_buf_1_im = r2Switch_10_out2_im;
  assign _zz_wn_re_3 = cnt_p1[8 : 0];
  assign _zz_wn_re_5 = _zz__zz_2_port0;
  assign _zz_wn_re_4 = _zz__zz_wn_re_4[23 : 0];
  assign _zz_wn_im_1 = _zz__zz_wn_im_1[23 : 0];
  assign r2Butterfly_11_wn_re = (mode ? _zz_wn_re_4 : _zz_wn_re_4);
  assign r2Butterfly_11_wn_im = (mode ? _zz_wn_im_1 : _zz_wn_im_12);
  assign r2Switch_11_sel = cnt[8];
  assign out0_buf_2_re = r2Switch_11_out1_re;
  assign out0_buf_2_im = r2Switch_11_out1_im;
  assign out1_buf_2_re = r2Switch_11_out2_re;
  assign out1_buf_2_im = r2Switch_11_out2_im;
  assign _zz_wn_re_6 = cnt_p1[7 : 0];
  assign _zz_wn_re_8 = _zz__zz_3_port0;
  assign _zz_wn_re_7 = _zz__zz_wn_re_7[23 : 0];
  assign _zz_wn_im_2 = _zz__zz_wn_im_2[23 : 0];
  assign r2Butterfly_12_wn_re = (mode ? _zz_wn_re_7 : _zz_wn_re_7);
  assign r2Butterfly_12_wn_im = (mode ? _zz_wn_im_2 : _zz_wn_im_14);
  assign r2Switch_12_sel = cnt[7];
  assign out0_buf_3_re = r2Switch_12_out1_re;
  assign out0_buf_3_im = r2Switch_12_out1_im;
  assign out1_buf_3_re = r2Switch_12_out2_re;
  assign out1_buf_3_im = r2Switch_12_out2_im;
  assign _zz_wn_re_9 = cnt_p1[6 : 0];
  assign _zz_wn_re_11 = _zz__zz_4_port0;
  assign _zz_wn_re_10 = _zz__zz_wn_re_10[23 : 0];
  assign _zz_wn_im_3 = _zz__zz_wn_im_3[23 : 0];
  assign r2Butterfly_13_wn_re = (mode ? _zz_wn_re_10 : _zz_wn_re_10);
  assign r2Butterfly_13_wn_im = (mode ? _zz_wn_im_3 : _zz_wn_im_16);
  assign r2Switch_13_sel = cnt[6];
  assign out0_buf_4_re = r2Switch_13_out1_re;
  assign out0_buf_4_im = r2Switch_13_out1_im;
  assign out1_buf_4_re = r2Switch_13_out2_re;
  assign out1_buf_4_im = r2Switch_13_out2_im;
  assign _zz_wn_re_12 = cnt_p1[5 : 0];
  assign _zz_wn_re_14 = _zz__zz_5_port0;
  assign _zz_wn_re_13 = _zz__zz_wn_re_13[23 : 0];
  assign _zz_wn_im_4 = _zz__zz_wn_im_4[23 : 0];
  assign r2Butterfly_14_wn_re = (mode ? _zz_wn_re_13 : _zz_wn_re_13);
  assign r2Butterfly_14_wn_im = (mode ? _zz_wn_im_4 : _zz_wn_im_18);
  assign r2Switch_14_sel = cnt[5];
  assign out0_buf_5_re = r2Switch_14_out1_re;
  assign out0_buf_5_im = r2Switch_14_out1_im;
  assign out1_buf_5_re = r2Switch_14_out2_re;
  assign out1_buf_5_im = r2Switch_14_out2_im;
  assign _zz_wn_re_15 = cnt_p1[4 : 0];
  assign _zz_wn_re_17 = _zz__zz_6_port0;
  assign _zz_wn_re_16 = _zz__zz_wn_re_16[23 : 0];
  assign _zz_wn_im_5 = _zz__zz_wn_im_5[23 : 0];
  assign r2Butterfly_15_wn_re = (mode ? _zz_wn_re_16 : _zz_wn_re_16);
  assign r2Butterfly_15_wn_im = (mode ? _zz_wn_im_5 : _zz_wn_im_20);
  assign r2Switch_15_sel = cnt[4];
  assign out0_buf_6_re = r2Switch_15_out1_re;
  assign out0_buf_6_im = r2Switch_15_out1_im;
  assign out1_buf_6_re = r2Switch_15_out2_re;
  assign out1_buf_6_im = r2Switch_15_out2_im;
  assign _zz_wn_re_18 = cnt_p1[3 : 0];
  assign _zz_wn_re_20 = _zz__zz_7_port0;
  assign _zz_wn_re_19 = _zz__zz_wn_re_19[23 : 0];
  assign _zz_wn_im_6 = _zz__zz_wn_im_6[23 : 0];
  assign r2Butterfly_16_wn_re = (mode ? _zz_wn_re_19 : _zz_wn_re_19);
  assign r2Butterfly_16_wn_im = (mode ? _zz_wn_im_6 : _zz_wn_im_22);
  assign r2Switch_16_sel = cnt[3];
  assign out0_buf_7_re = r2Switch_16_out1_re;
  assign out0_buf_7_im = r2Switch_16_out1_im;
  assign out1_buf_7_re = r2Switch_16_out2_re;
  assign out1_buf_7_im = r2Switch_16_out2_im;
  assign _zz_wn_re_21 = cnt_p1[2 : 0];
  assign _zz_wn_re_23 = _zz__zz_8_port0;
  assign _zz_wn_re_22 = _zz__zz_wn_re_22[23 : 0];
  assign _zz_wn_im_7 = _zz__zz_wn_im_7[23 : 0];
  assign r2Butterfly_17_wn_re = (mode ? _zz_wn_re_22 : _zz_wn_re_22);
  assign r2Butterfly_17_wn_im = (mode ? _zz_wn_im_7 : _zz_wn_im_24);
  assign r2Switch_17_sel = cnt[2];
  assign out0_buf_8_re = r2Switch_17_out1_re;
  assign out0_buf_8_im = r2Switch_17_out1_im;
  assign out1_buf_8_re = r2Switch_17_out2_re;
  assign out1_buf_8_im = r2Switch_17_out2_im;
  assign _zz_wn_re_24 = cnt_p1[1 : 0];
  assign _zz_wn_re_26 = _zz__zz_9_port0;
  assign _zz_wn_re_25 = _zz__zz_wn_re_25[23 : 0];
  assign _zz_wn_im_8 = _zz__zz_wn_im_8[23 : 0];
  assign r2Butterfly_18_wn_re = (mode ? _zz_wn_re_25 : _zz_wn_re_25);
  assign r2Butterfly_18_wn_im = (mode ? _zz_wn_im_8 : _zz_wn_im_26);
  assign r2Switch_18_sel = cnt[1];
  assign out0_buf_9_re = r2Switch_18_out1_re;
  assign out0_buf_9_im = r2Switch_18_out1_im;
  assign out1_buf_9_re = r2Switch_18_out2_re;
  assign out1_buf_9_im = r2Switch_18_out2_im;
  assign _zz_wn_re_27 = cnt_p1[0 : 0];
  assign _zz_wn_re_29 = _zz__zz_10_port0;
  assign _zz_wn_re_28 = _zz__zz_wn_re_28[23 : 0];
  assign _zz_wn_im_9 = _zz__zz_wn_im_9[23 : 0];
  assign r2Butterfly_19_wn_re = (mode ? _zz_wn_re_28 : _zz_wn_re_28);
  assign r2Butterfly_19_wn_im = (mode ? _zz_wn_im_9 : _zz_wn_im_28);
  assign r2Switch_19_sel = cnt[0];
  assign out0_buf_10_re = r2Switch_19_out1_re;
  assign out0_buf_10_im = r2Switch_19_out1_im;
  assign out1_buf_10_re = r2Switch_19_out2_re;
  assign out1_buf_10_im = r2Switch_19_out2_im;
  assign out0_buf_11_re = ($signed(out1D1_re) + $signed(out1_buf_10_re));
  assign out0_buf_11_im = ($signed(out1D1_im) + $signed(out1_buf_10_im));
  assign out1_buf_11_re = ($signed(out1D1_re) - $signed(out1_buf_10_re));
  assign out1_buf_11_im = ($signed(out1D1_im) - $signed(out1_buf_10_im));
  assign result_out1_re = (mode ? out0_buf_11_re : _zz_result_out1_re);
  assign result_out1_im = (mode ? out0_buf_11_im : _zz_result_out1_im);
  assign result_out2_re = (mode ? out1_buf_11_re : _zz_result_out2_re);
  assign result_out2_im = (mode ? out1_buf_11_im : _zz_result_out2_im);
  assign reorder_1_unsorted_valid = (12'h7ff < cnt);
  assign result_valid = reorder_1_sorted_valid;
  assign result_payload_last = reorder_1_sorted_payload_last;
  assign result_payload_fragment_re = reorder_1_sorted_payload_fragment_re;
  assign result_payload_fragment_im = reorder_1_sorted_payload_fragment_im;
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      cnt <= 12'h0;
    end else begin
      if(when_R2MDC_l20) begin
        cnt <= ((cnt == 12'hbff) ? 12'h0 : _zz_cnt);
      end
    end
  end

  always @(posedge clk) begin
    out1D1_re <= out0_buf_10_re;
    out1D1_im <= out0_buf_10_im;
    result_out1_regNext_re <= result_out1_re;
    result_out1_regNext_im <= result_out1_im;
    result_out2_regNext_re <= result_out2_re;
    result_out2_regNext_im <= result_out2_im;
  end


endmodule

module Reorder (
  input               unsorted_valid,
  input      [23:0]   unsorted_payload_in0_re,
  input      [23:0]   unsorted_payload_in0_im,
  input      [23:0]   unsorted_payload_in1_re,
  input      [23:0]   unsorted_payload_in1_im,
  output              sorted_valid,
  output              sorted_payload_last,
  output reg [23:0]   sorted_payload_fragment_re,
  output reg [23:0]   sorted_payload_fragment_im,
  input               clk,
  input               reset
);
  reg        [47:0]   _zz_ram_low_port1;
  reg        [47:0]   _zz_ram_high_port1;
  wire       [47:0]   _zz_ram_low_port;
  wire       [47:0]   _zz_ram_high_port;
  wire       [9:0]    _zz__zz_sorted_payload_fragment_re_1;
  wire                _zz__zz_sorted_payload_fragment_re_1_1;
  wire       [23:0]   _zz_sorted_payload_fragment_re_4;
  wire       [23:0]   _zz_sorted_payload_fragment_im;
  wire       [9:0]    _zz__zz_sorted_payload_fragment_re_3;
  wire                _zz__zz_sorted_payload_fragment_re_3_1;
  wire       [23:0]   _zz_sorted_payload_fragment_re_5;
  wire       [23:0]   _zz_sorted_payload_fragment_im_1;
  wire       [9:0]    _zz_ram_low_port_1;
  wire                _zz_ram_low_port_2;
  wire       [9:0]    _zz_ram_high_port_1;
  wire                _zz_ram_high_port_2;
  reg                 _zz_1;
  reg                 _zz_2;
  reg        [9:0]    in_cnt;
  reg        [10:0]   out_cnt;
  wire       [9:0]    in_cnt_index;
  wire                sorted_valid_1;
  reg                 _zz_3;
  wire       [10:0]   _zz_sorted_payload_fragment_re;
  wire       [47:0]   _zz_sorted_payload_fragment_re_1;
  wire       [10:0]   _zz_sorted_payload_fragment_re_2;
  wire       [47:0]   _zz_sorted_payload_fragment_re_3;
  reg                 sorted_valid_1_regNext;
  (* ram_style = "block" *) reg [47:0] ram_low [0:1023];
  (* ram_style = "block" *) reg [47:0] ram_high [0:1023];

  assign _zz_ram_low_port_1 = _zz_sorted_payload_fragment_re[9:0];
  assign _zz_sorted_payload_fragment_re_4 = _zz_sorted_payload_fragment_re_1[23 : 0];
  assign _zz_sorted_payload_fragment_im = _zz_sorted_payload_fragment_re_1[47 : 24];
  assign _zz_ram_high_port_1 = _zz_sorted_payload_fragment_re_2[9:0];
  assign _zz_sorted_payload_fragment_re_5 = _zz_sorted_payload_fragment_re_3[23 : 0];
  assign _zz_sorted_payload_fragment_im_1 = _zz_sorted_payload_fragment_re_3[47 : 24];
  assign _zz_ram_low_port = {unsorted_payload_in0_im,unsorted_payload_in0_re};
  assign _zz_ram_low_port_2 = 1'b1;
  assign _zz_ram_high_port = {unsorted_payload_in1_im,unsorted_payload_in1_re};
  assign _zz_ram_high_port_2 = 1'b1;
  always @(posedge clk) begin
    if(_zz_2) begin
      ram_low[in_cnt_index] <= _zz_ram_low_port;
    end
  end

  always @(posedge clk) begin
    if(_zz_ram_low_port_2) begin
      _zz_ram_low_port1 <= ram_low[_zz_ram_low_port_1];
    end
  end

  always @(posedge clk) begin
    if(_zz_1) begin
      ram_high[in_cnt_index] <= _zz_ram_high_port;
    end
  end

  always @(posedge clk) begin
    if(_zz_ram_high_port_2) begin
      _zz_ram_high_port1 <= ram_high[_zz_ram_high_port_1];
    end
  end

  always @(*) begin
    _zz_1 = 1'b0;
    if(unsorted_valid) begin
      _zz_1 = 1'b1;
    end
  end

  always @(*) begin
    _zz_2 = 1'b0;
    if(unsorted_valid) begin
      _zz_2 = 1'b1;
    end
  end

  assign in_cnt_index = {in_cnt[0],{in_cnt[1],{in_cnt[2],{in_cnt[3],{in_cnt[4],{in_cnt[5],{in_cnt[6],{in_cnt[7],{in_cnt[8],in_cnt[9]}}}}}}}}};
  assign sorted_valid_1 = ((in_cnt == 10'h3ff) || (out_cnt != 11'h0));
  assign _zz_sorted_payload_fragment_re = out_cnt;
  assign _zz_sorted_payload_fragment_re_1 = _zz_ram_low_port1;
  always @(*) begin
    if(_zz_3) begin
      sorted_payload_fragment_re = _zz_sorted_payload_fragment_re_4[23 : 0];
    end else begin
      sorted_payload_fragment_re = _zz_sorted_payload_fragment_re_5[23 : 0];
    end
  end

  always @(*) begin
    if(_zz_3) begin
      sorted_payload_fragment_im = _zz_sorted_payload_fragment_im[23 : 0];
    end else begin
      sorted_payload_fragment_im = _zz_sorted_payload_fragment_im_1[23 : 0];
    end
  end

  assign _zz_sorted_payload_fragment_re_2 = out_cnt;
  assign _zz_sorted_payload_fragment_re_3 = _zz_ram_high_port1;
  assign sorted_payload_last = ((out_cnt == 11'h0) && sorted_valid);
  assign sorted_valid = sorted_valid_1_regNext;
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      in_cnt <= 10'h0;
      out_cnt <= 11'h0;
    end else begin
      if(unsorted_valid) begin
        in_cnt <= (in_cnt + 10'h001);
      end
      if(sorted_valid_1) begin
        out_cnt <= (out_cnt + 11'h001);
      end
    end
  end

  always @(posedge clk) begin
    _zz_3 <= (out_cnt < 11'h400);
    sorted_valid_1_regNext <= sorted_valid_1;
  end


endmodule

//R2Switch replaced by R2Switch

module ShiftRegisterNE_19 (
  input      [23:0]   input_re,
  input      [23:0]   input_im,
  output     [23:0]   output_re,
  output     [23:0]   output_im,
  input               clk,
  input               reset
);
  reg        [23:0]   shift_reg_0_re;
  reg        [23:0]   shift_reg_0_im;

  assign output_re = shift_reg_0_re;
  assign output_im = shift_reg_0_im;
  always @(posedge clk) begin
    shift_reg_0_re <= input_re;
    shift_reg_0_im <= input_im;
  end


endmodule

//R2Butterfly replaced by R2Butterfly

//ShiftRegisterNE_17 replaced by ShiftRegisterNE_17

//R2Switch replaced by R2Switch

module ShiftRegisterNE_17 (
  input      [23:0]   input_re,
  input      [23:0]   input_im,
  output     [23:0]   output_re,
  output     [23:0]   output_im,
  input               clk,
  input               reset
);
  reg        [23:0]   shift_reg_0_re;
  reg        [23:0]   shift_reg_0_im;
  reg        [23:0]   shift_reg_1_re;
  reg        [23:0]   shift_reg_1_im;

  assign output_re = shift_reg_1_re;
  assign output_im = shift_reg_1_im;
  always @(posedge clk) begin
    shift_reg_0_re <= input_re;
    shift_reg_0_im <= input_im;
    shift_reg_1_re <= shift_reg_0_re;
    shift_reg_1_im <= shift_reg_0_im;
  end


endmodule

//R2Butterfly replaced by R2Butterfly

//ShiftRegisterNE_15 replaced by ShiftRegisterNE_15

//R2Switch replaced by R2Switch

module ShiftRegisterNE_15 (
  input      [23:0]   input_re,
  input      [23:0]   input_im,
  output     [23:0]   output_re,
  output     [23:0]   output_im,
  input               clk,
  input               reset
);
  reg        [23:0]   shift_reg_0_re;
  reg        [23:0]   shift_reg_0_im;
  reg        [23:0]   shift_reg_1_re;
  reg        [23:0]   shift_reg_1_im;
  reg        [23:0]   shift_reg_2_re;
  reg        [23:0]   shift_reg_2_im;
  reg        [23:0]   shift_reg_3_re;
  reg        [23:0]   shift_reg_3_im;

  assign output_re = shift_reg_3_re;
  assign output_im = shift_reg_3_im;
  always @(posedge clk) begin
    shift_reg_0_re <= input_re;
    shift_reg_0_im <= input_im;
    shift_reg_1_re <= shift_reg_0_re;
    shift_reg_1_im <= shift_reg_0_im;
    shift_reg_2_re <= shift_reg_1_re;
    shift_reg_2_im <= shift_reg_1_im;
    shift_reg_3_re <= shift_reg_2_re;
    shift_reg_3_im <= shift_reg_2_im;
  end


endmodule

//R2Butterfly replaced by R2Butterfly

//ShiftRegisterNE_13 replaced by ShiftRegisterNE_13

//R2Switch replaced by R2Switch

module ShiftRegisterNE_13 (
  input      [23:0]   input_re,
  input      [23:0]   input_im,
  output     [23:0]   output_re,
  output     [23:0]   output_im,
  input               clk,
  input               reset
);
  reg        [23:0]   shift_reg_0_re;
  reg        [23:0]   shift_reg_0_im;
  reg        [23:0]   shift_reg_1_re;
  reg        [23:0]   shift_reg_1_im;
  reg        [23:0]   shift_reg_2_re;
  reg        [23:0]   shift_reg_2_im;
  reg        [23:0]   shift_reg_3_re;
  reg        [23:0]   shift_reg_3_im;
  reg        [23:0]   shift_reg_4_re;
  reg        [23:0]   shift_reg_4_im;
  reg        [23:0]   shift_reg_5_re;
  reg        [23:0]   shift_reg_5_im;
  reg        [23:0]   shift_reg_6_re;
  reg        [23:0]   shift_reg_6_im;
  reg        [23:0]   shift_reg_7_re;
  reg        [23:0]   shift_reg_7_im;

  assign output_re = shift_reg_7_re;
  assign output_im = shift_reg_7_im;
  always @(posedge clk) begin
    shift_reg_0_re <= input_re;
    shift_reg_0_im <= input_im;
    shift_reg_1_re <= shift_reg_0_re;
    shift_reg_1_im <= shift_reg_0_im;
    shift_reg_2_re <= shift_reg_1_re;
    shift_reg_2_im <= shift_reg_1_im;
    shift_reg_3_re <= shift_reg_2_re;
    shift_reg_3_im <= shift_reg_2_im;
    shift_reg_4_re <= shift_reg_3_re;
    shift_reg_4_im <= shift_reg_3_im;
    shift_reg_5_re <= shift_reg_4_re;
    shift_reg_5_im <= shift_reg_4_im;
    shift_reg_6_re <= shift_reg_5_re;
    shift_reg_6_im <= shift_reg_5_im;
    shift_reg_7_re <= shift_reg_6_re;
    shift_reg_7_im <= shift_reg_6_im;
  end


endmodule

//R2Butterfly replaced by R2Butterfly

//ShiftRegisterNE_11 replaced by ShiftRegisterNE_11

//R2Switch replaced by R2Switch

module ShiftRegisterNE_11 (
  input      [23:0]   input_re,
  input      [23:0]   input_im,
  output     [23:0]   output_re,
  output     [23:0]   output_im,
  input               clk,
  input               reset
);
  reg        [23:0]   shift_reg_0_re;
  reg        [23:0]   shift_reg_0_im;
  reg        [23:0]   shift_reg_1_re;
  reg        [23:0]   shift_reg_1_im;
  reg        [23:0]   shift_reg_2_re;
  reg        [23:0]   shift_reg_2_im;
  reg        [23:0]   shift_reg_3_re;
  reg        [23:0]   shift_reg_3_im;
  reg        [23:0]   shift_reg_4_re;
  reg        [23:0]   shift_reg_4_im;
  reg        [23:0]   shift_reg_5_re;
  reg        [23:0]   shift_reg_5_im;
  reg        [23:0]   shift_reg_6_re;
  reg        [23:0]   shift_reg_6_im;
  reg        [23:0]   shift_reg_7_re;
  reg        [23:0]   shift_reg_7_im;
  reg        [23:0]   shift_reg_8_re;
  reg        [23:0]   shift_reg_8_im;
  reg        [23:0]   shift_reg_9_re;
  reg        [23:0]   shift_reg_9_im;
  reg        [23:0]   shift_reg_10_re;
  reg        [23:0]   shift_reg_10_im;
  reg        [23:0]   shift_reg_11_re;
  reg        [23:0]   shift_reg_11_im;
  reg        [23:0]   shift_reg_12_re;
  reg        [23:0]   shift_reg_12_im;
  reg        [23:0]   shift_reg_13_re;
  reg        [23:0]   shift_reg_13_im;
  reg        [23:0]   shift_reg_14_re;
  reg        [23:0]   shift_reg_14_im;
  reg        [23:0]   shift_reg_15_re;
  reg        [23:0]   shift_reg_15_im;

  assign output_re = shift_reg_15_re;
  assign output_im = shift_reg_15_im;
  always @(posedge clk) begin
    shift_reg_0_re <= input_re;
    shift_reg_0_im <= input_im;
    shift_reg_1_re <= shift_reg_0_re;
    shift_reg_1_im <= shift_reg_0_im;
    shift_reg_2_re <= shift_reg_1_re;
    shift_reg_2_im <= shift_reg_1_im;
    shift_reg_3_re <= shift_reg_2_re;
    shift_reg_3_im <= shift_reg_2_im;
    shift_reg_4_re <= shift_reg_3_re;
    shift_reg_4_im <= shift_reg_3_im;
    shift_reg_5_re <= shift_reg_4_re;
    shift_reg_5_im <= shift_reg_4_im;
    shift_reg_6_re <= shift_reg_5_re;
    shift_reg_6_im <= shift_reg_5_im;
    shift_reg_7_re <= shift_reg_6_re;
    shift_reg_7_im <= shift_reg_6_im;
    shift_reg_8_re <= shift_reg_7_re;
    shift_reg_8_im <= shift_reg_7_im;
    shift_reg_9_re <= shift_reg_8_re;
    shift_reg_9_im <= shift_reg_8_im;
    shift_reg_10_re <= shift_reg_9_re;
    shift_reg_10_im <= shift_reg_9_im;
    shift_reg_11_re <= shift_reg_10_re;
    shift_reg_11_im <= shift_reg_10_im;
    shift_reg_12_re <= shift_reg_11_re;
    shift_reg_12_im <= shift_reg_11_im;
    shift_reg_13_re <= shift_reg_12_re;
    shift_reg_13_im <= shift_reg_12_im;
    shift_reg_14_re <= shift_reg_13_re;
    shift_reg_14_im <= shift_reg_13_im;
    shift_reg_15_re <= shift_reg_14_re;
    shift_reg_15_im <= shift_reg_14_im;
  end


endmodule

//R2Butterfly replaced by R2Butterfly

//ShiftRegisterNE_9 replaced by ShiftRegisterNE_9

//R2Switch replaced by R2Switch

module ShiftRegisterNE_9 (
  input      [23:0]   input_re,
  input      [23:0]   input_im,
  output     [23:0]   output_re,
  output     [23:0]   output_im,
  input               clk,
  input               reset
);
  reg        [23:0]   shift_reg_0_re;
  reg        [23:0]   shift_reg_0_im;
  reg        [23:0]   shift_reg_1_re;
  reg        [23:0]   shift_reg_1_im;
  reg        [23:0]   shift_reg_2_re;
  reg        [23:0]   shift_reg_2_im;
  reg        [23:0]   shift_reg_3_re;
  reg        [23:0]   shift_reg_3_im;
  reg        [23:0]   shift_reg_4_re;
  reg        [23:0]   shift_reg_4_im;
  reg        [23:0]   shift_reg_5_re;
  reg        [23:0]   shift_reg_5_im;
  reg        [23:0]   shift_reg_6_re;
  reg        [23:0]   shift_reg_6_im;
  reg        [23:0]   shift_reg_7_re;
  reg        [23:0]   shift_reg_7_im;
  reg        [23:0]   shift_reg_8_re;
  reg        [23:0]   shift_reg_8_im;
  reg        [23:0]   shift_reg_9_re;
  reg        [23:0]   shift_reg_9_im;
  reg        [23:0]   shift_reg_10_re;
  reg        [23:0]   shift_reg_10_im;
  reg        [23:0]   shift_reg_11_re;
  reg        [23:0]   shift_reg_11_im;
  reg        [23:0]   shift_reg_12_re;
  reg        [23:0]   shift_reg_12_im;
  reg        [23:0]   shift_reg_13_re;
  reg        [23:0]   shift_reg_13_im;
  reg        [23:0]   shift_reg_14_re;
  reg        [23:0]   shift_reg_14_im;
  reg        [23:0]   shift_reg_15_re;
  reg        [23:0]   shift_reg_15_im;
  reg        [23:0]   shift_reg_16_re;
  reg        [23:0]   shift_reg_16_im;
  reg        [23:0]   shift_reg_17_re;
  reg        [23:0]   shift_reg_17_im;
  reg        [23:0]   shift_reg_18_re;
  reg        [23:0]   shift_reg_18_im;
  reg        [23:0]   shift_reg_19_re;
  reg        [23:0]   shift_reg_19_im;
  reg        [23:0]   shift_reg_20_re;
  reg        [23:0]   shift_reg_20_im;
  reg        [23:0]   shift_reg_21_re;
  reg        [23:0]   shift_reg_21_im;
  reg        [23:0]   shift_reg_22_re;
  reg        [23:0]   shift_reg_22_im;
  reg        [23:0]   shift_reg_23_re;
  reg        [23:0]   shift_reg_23_im;
  reg        [23:0]   shift_reg_24_re;
  reg        [23:0]   shift_reg_24_im;
  reg        [23:0]   shift_reg_25_re;
  reg        [23:0]   shift_reg_25_im;
  reg        [23:0]   shift_reg_26_re;
  reg        [23:0]   shift_reg_26_im;
  reg        [23:0]   shift_reg_27_re;
  reg        [23:0]   shift_reg_27_im;
  reg        [23:0]   shift_reg_28_re;
  reg        [23:0]   shift_reg_28_im;
  reg        [23:0]   shift_reg_29_re;
  reg        [23:0]   shift_reg_29_im;
  reg        [23:0]   shift_reg_30_re;
  reg        [23:0]   shift_reg_30_im;
  reg        [23:0]   shift_reg_31_re;
  reg        [23:0]   shift_reg_31_im;

  assign output_re = shift_reg_31_re;
  assign output_im = shift_reg_31_im;
  always @(posedge clk) begin
    shift_reg_0_re <= input_re;
    shift_reg_0_im <= input_im;
    shift_reg_1_re <= shift_reg_0_re;
    shift_reg_1_im <= shift_reg_0_im;
    shift_reg_2_re <= shift_reg_1_re;
    shift_reg_2_im <= shift_reg_1_im;
    shift_reg_3_re <= shift_reg_2_re;
    shift_reg_3_im <= shift_reg_2_im;
    shift_reg_4_re <= shift_reg_3_re;
    shift_reg_4_im <= shift_reg_3_im;
    shift_reg_5_re <= shift_reg_4_re;
    shift_reg_5_im <= shift_reg_4_im;
    shift_reg_6_re <= shift_reg_5_re;
    shift_reg_6_im <= shift_reg_5_im;
    shift_reg_7_re <= shift_reg_6_re;
    shift_reg_7_im <= shift_reg_6_im;
    shift_reg_8_re <= shift_reg_7_re;
    shift_reg_8_im <= shift_reg_7_im;
    shift_reg_9_re <= shift_reg_8_re;
    shift_reg_9_im <= shift_reg_8_im;
    shift_reg_10_re <= shift_reg_9_re;
    shift_reg_10_im <= shift_reg_9_im;
    shift_reg_11_re <= shift_reg_10_re;
    shift_reg_11_im <= shift_reg_10_im;
    shift_reg_12_re <= shift_reg_11_re;
    shift_reg_12_im <= shift_reg_11_im;
    shift_reg_13_re <= shift_reg_12_re;
    shift_reg_13_im <= shift_reg_12_im;
    shift_reg_14_re <= shift_reg_13_re;
    shift_reg_14_im <= shift_reg_13_im;
    shift_reg_15_re <= shift_reg_14_re;
    shift_reg_15_im <= shift_reg_14_im;
    shift_reg_16_re <= shift_reg_15_re;
    shift_reg_16_im <= shift_reg_15_im;
    shift_reg_17_re <= shift_reg_16_re;
    shift_reg_17_im <= shift_reg_16_im;
    shift_reg_18_re <= shift_reg_17_re;
    shift_reg_18_im <= shift_reg_17_im;
    shift_reg_19_re <= shift_reg_18_re;
    shift_reg_19_im <= shift_reg_18_im;
    shift_reg_20_re <= shift_reg_19_re;
    shift_reg_20_im <= shift_reg_19_im;
    shift_reg_21_re <= shift_reg_20_re;
    shift_reg_21_im <= shift_reg_20_im;
    shift_reg_22_re <= shift_reg_21_re;
    shift_reg_22_im <= shift_reg_21_im;
    shift_reg_23_re <= shift_reg_22_re;
    shift_reg_23_im <= shift_reg_22_im;
    shift_reg_24_re <= shift_reg_23_re;
    shift_reg_24_im <= shift_reg_23_im;
    shift_reg_25_re <= shift_reg_24_re;
    shift_reg_25_im <= shift_reg_24_im;
    shift_reg_26_re <= shift_reg_25_re;
    shift_reg_26_im <= shift_reg_25_im;
    shift_reg_27_re <= shift_reg_26_re;
    shift_reg_27_im <= shift_reg_26_im;
    shift_reg_28_re <= shift_reg_27_re;
    shift_reg_28_im <= shift_reg_27_im;
    shift_reg_29_re <= shift_reg_28_re;
    shift_reg_29_im <= shift_reg_28_im;
    shift_reg_30_re <= shift_reg_29_re;
    shift_reg_30_im <= shift_reg_29_im;
    shift_reg_31_re <= shift_reg_30_re;
    shift_reg_31_im <= shift_reg_30_im;
  end


endmodule

//R2Butterfly replaced by R2Butterfly

//ShiftRegisterNE_7 replaced by ShiftRegisterNE_7

//R2Switch replaced by R2Switch

module ShiftRegisterNE_7 (
  input      [23:0]   input_re,
  input      [23:0]   input_im,
  output     [23:0]   output_re,
  output     [23:0]   output_im,
  input               clk,
  input               reset
);
  reg        [23:0]   shift_reg_0_re;
  reg        [23:0]   shift_reg_0_im;
  reg        [23:0]   shift_reg_1_re;
  reg        [23:0]   shift_reg_1_im;
  reg        [23:0]   shift_reg_2_re;
  reg        [23:0]   shift_reg_2_im;
  reg        [23:0]   shift_reg_3_re;
  reg        [23:0]   shift_reg_3_im;
  reg        [23:0]   shift_reg_4_re;
  reg        [23:0]   shift_reg_4_im;
  reg        [23:0]   shift_reg_5_re;
  reg        [23:0]   shift_reg_5_im;
  reg        [23:0]   shift_reg_6_re;
  reg        [23:0]   shift_reg_6_im;
  reg        [23:0]   shift_reg_7_re;
  reg        [23:0]   shift_reg_7_im;
  reg        [23:0]   shift_reg_8_re;
  reg        [23:0]   shift_reg_8_im;
  reg        [23:0]   shift_reg_9_re;
  reg        [23:0]   shift_reg_9_im;
  reg        [23:0]   shift_reg_10_re;
  reg        [23:0]   shift_reg_10_im;
  reg        [23:0]   shift_reg_11_re;
  reg        [23:0]   shift_reg_11_im;
  reg        [23:0]   shift_reg_12_re;
  reg        [23:0]   shift_reg_12_im;
  reg        [23:0]   shift_reg_13_re;
  reg        [23:0]   shift_reg_13_im;
  reg        [23:0]   shift_reg_14_re;
  reg        [23:0]   shift_reg_14_im;
  reg        [23:0]   shift_reg_15_re;
  reg        [23:0]   shift_reg_15_im;
  reg        [23:0]   shift_reg_16_re;
  reg        [23:0]   shift_reg_16_im;
  reg        [23:0]   shift_reg_17_re;
  reg        [23:0]   shift_reg_17_im;
  reg        [23:0]   shift_reg_18_re;
  reg        [23:0]   shift_reg_18_im;
  reg        [23:0]   shift_reg_19_re;
  reg        [23:0]   shift_reg_19_im;
  reg        [23:0]   shift_reg_20_re;
  reg        [23:0]   shift_reg_20_im;
  reg        [23:0]   shift_reg_21_re;
  reg        [23:0]   shift_reg_21_im;
  reg        [23:0]   shift_reg_22_re;
  reg        [23:0]   shift_reg_22_im;
  reg        [23:0]   shift_reg_23_re;
  reg        [23:0]   shift_reg_23_im;
  reg        [23:0]   shift_reg_24_re;
  reg        [23:0]   shift_reg_24_im;
  reg        [23:0]   shift_reg_25_re;
  reg        [23:0]   shift_reg_25_im;
  reg        [23:0]   shift_reg_26_re;
  reg        [23:0]   shift_reg_26_im;
  reg        [23:0]   shift_reg_27_re;
  reg        [23:0]   shift_reg_27_im;
  reg        [23:0]   shift_reg_28_re;
  reg        [23:0]   shift_reg_28_im;
  reg        [23:0]   shift_reg_29_re;
  reg        [23:0]   shift_reg_29_im;
  reg        [23:0]   shift_reg_30_re;
  reg        [23:0]   shift_reg_30_im;
  reg        [23:0]   shift_reg_31_re;
  reg        [23:0]   shift_reg_31_im;
  reg        [23:0]   shift_reg_32_re;
  reg        [23:0]   shift_reg_32_im;
  reg        [23:0]   shift_reg_33_re;
  reg        [23:0]   shift_reg_33_im;
  reg        [23:0]   shift_reg_34_re;
  reg        [23:0]   shift_reg_34_im;
  reg        [23:0]   shift_reg_35_re;
  reg        [23:0]   shift_reg_35_im;
  reg        [23:0]   shift_reg_36_re;
  reg        [23:0]   shift_reg_36_im;
  reg        [23:0]   shift_reg_37_re;
  reg        [23:0]   shift_reg_37_im;
  reg        [23:0]   shift_reg_38_re;
  reg        [23:0]   shift_reg_38_im;
  reg        [23:0]   shift_reg_39_re;
  reg        [23:0]   shift_reg_39_im;
  reg        [23:0]   shift_reg_40_re;
  reg        [23:0]   shift_reg_40_im;
  reg        [23:0]   shift_reg_41_re;
  reg        [23:0]   shift_reg_41_im;
  reg        [23:0]   shift_reg_42_re;
  reg        [23:0]   shift_reg_42_im;
  reg        [23:0]   shift_reg_43_re;
  reg        [23:0]   shift_reg_43_im;
  reg        [23:0]   shift_reg_44_re;
  reg        [23:0]   shift_reg_44_im;
  reg        [23:0]   shift_reg_45_re;
  reg        [23:0]   shift_reg_45_im;
  reg        [23:0]   shift_reg_46_re;
  reg        [23:0]   shift_reg_46_im;
  reg        [23:0]   shift_reg_47_re;
  reg        [23:0]   shift_reg_47_im;
  reg        [23:0]   shift_reg_48_re;
  reg        [23:0]   shift_reg_48_im;
  reg        [23:0]   shift_reg_49_re;
  reg        [23:0]   shift_reg_49_im;
  reg        [23:0]   shift_reg_50_re;
  reg        [23:0]   shift_reg_50_im;
  reg        [23:0]   shift_reg_51_re;
  reg        [23:0]   shift_reg_51_im;
  reg        [23:0]   shift_reg_52_re;
  reg        [23:0]   shift_reg_52_im;
  reg        [23:0]   shift_reg_53_re;
  reg        [23:0]   shift_reg_53_im;
  reg        [23:0]   shift_reg_54_re;
  reg        [23:0]   shift_reg_54_im;
  reg        [23:0]   shift_reg_55_re;
  reg        [23:0]   shift_reg_55_im;
  reg        [23:0]   shift_reg_56_re;
  reg        [23:0]   shift_reg_56_im;
  reg        [23:0]   shift_reg_57_re;
  reg        [23:0]   shift_reg_57_im;
  reg        [23:0]   shift_reg_58_re;
  reg        [23:0]   shift_reg_58_im;
  reg        [23:0]   shift_reg_59_re;
  reg        [23:0]   shift_reg_59_im;
  reg        [23:0]   shift_reg_60_re;
  reg        [23:0]   shift_reg_60_im;
  reg        [23:0]   shift_reg_61_re;
  reg        [23:0]   shift_reg_61_im;
  reg        [23:0]   shift_reg_62_re;
  reg        [23:0]   shift_reg_62_im;
  reg        [23:0]   shift_reg_63_re;
  reg        [23:0]   shift_reg_63_im;

  assign output_re = shift_reg_63_re;
  assign output_im = shift_reg_63_im;
  always @(posedge clk) begin
    shift_reg_0_re <= input_re;
    shift_reg_0_im <= input_im;
    shift_reg_1_re <= shift_reg_0_re;
    shift_reg_1_im <= shift_reg_0_im;
    shift_reg_2_re <= shift_reg_1_re;
    shift_reg_2_im <= shift_reg_1_im;
    shift_reg_3_re <= shift_reg_2_re;
    shift_reg_3_im <= shift_reg_2_im;
    shift_reg_4_re <= shift_reg_3_re;
    shift_reg_4_im <= shift_reg_3_im;
    shift_reg_5_re <= shift_reg_4_re;
    shift_reg_5_im <= shift_reg_4_im;
    shift_reg_6_re <= shift_reg_5_re;
    shift_reg_6_im <= shift_reg_5_im;
    shift_reg_7_re <= shift_reg_6_re;
    shift_reg_7_im <= shift_reg_6_im;
    shift_reg_8_re <= shift_reg_7_re;
    shift_reg_8_im <= shift_reg_7_im;
    shift_reg_9_re <= shift_reg_8_re;
    shift_reg_9_im <= shift_reg_8_im;
    shift_reg_10_re <= shift_reg_9_re;
    shift_reg_10_im <= shift_reg_9_im;
    shift_reg_11_re <= shift_reg_10_re;
    shift_reg_11_im <= shift_reg_10_im;
    shift_reg_12_re <= shift_reg_11_re;
    shift_reg_12_im <= shift_reg_11_im;
    shift_reg_13_re <= shift_reg_12_re;
    shift_reg_13_im <= shift_reg_12_im;
    shift_reg_14_re <= shift_reg_13_re;
    shift_reg_14_im <= shift_reg_13_im;
    shift_reg_15_re <= shift_reg_14_re;
    shift_reg_15_im <= shift_reg_14_im;
    shift_reg_16_re <= shift_reg_15_re;
    shift_reg_16_im <= shift_reg_15_im;
    shift_reg_17_re <= shift_reg_16_re;
    shift_reg_17_im <= shift_reg_16_im;
    shift_reg_18_re <= shift_reg_17_re;
    shift_reg_18_im <= shift_reg_17_im;
    shift_reg_19_re <= shift_reg_18_re;
    shift_reg_19_im <= shift_reg_18_im;
    shift_reg_20_re <= shift_reg_19_re;
    shift_reg_20_im <= shift_reg_19_im;
    shift_reg_21_re <= shift_reg_20_re;
    shift_reg_21_im <= shift_reg_20_im;
    shift_reg_22_re <= shift_reg_21_re;
    shift_reg_22_im <= shift_reg_21_im;
    shift_reg_23_re <= shift_reg_22_re;
    shift_reg_23_im <= shift_reg_22_im;
    shift_reg_24_re <= shift_reg_23_re;
    shift_reg_24_im <= shift_reg_23_im;
    shift_reg_25_re <= shift_reg_24_re;
    shift_reg_25_im <= shift_reg_24_im;
    shift_reg_26_re <= shift_reg_25_re;
    shift_reg_26_im <= shift_reg_25_im;
    shift_reg_27_re <= shift_reg_26_re;
    shift_reg_27_im <= shift_reg_26_im;
    shift_reg_28_re <= shift_reg_27_re;
    shift_reg_28_im <= shift_reg_27_im;
    shift_reg_29_re <= shift_reg_28_re;
    shift_reg_29_im <= shift_reg_28_im;
    shift_reg_30_re <= shift_reg_29_re;
    shift_reg_30_im <= shift_reg_29_im;
    shift_reg_31_re <= shift_reg_30_re;
    shift_reg_31_im <= shift_reg_30_im;
    shift_reg_32_re <= shift_reg_31_re;
    shift_reg_32_im <= shift_reg_31_im;
    shift_reg_33_re <= shift_reg_32_re;
    shift_reg_33_im <= shift_reg_32_im;
    shift_reg_34_re <= shift_reg_33_re;
    shift_reg_34_im <= shift_reg_33_im;
    shift_reg_35_re <= shift_reg_34_re;
    shift_reg_35_im <= shift_reg_34_im;
    shift_reg_36_re <= shift_reg_35_re;
    shift_reg_36_im <= shift_reg_35_im;
    shift_reg_37_re <= shift_reg_36_re;
    shift_reg_37_im <= shift_reg_36_im;
    shift_reg_38_re <= shift_reg_37_re;
    shift_reg_38_im <= shift_reg_37_im;
    shift_reg_39_re <= shift_reg_38_re;
    shift_reg_39_im <= shift_reg_38_im;
    shift_reg_40_re <= shift_reg_39_re;
    shift_reg_40_im <= shift_reg_39_im;
    shift_reg_41_re <= shift_reg_40_re;
    shift_reg_41_im <= shift_reg_40_im;
    shift_reg_42_re <= shift_reg_41_re;
    shift_reg_42_im <= shift_reg_41_im;
    shift_reg_43_re <= shift_reg_42_re;
    shift_reg_43_im <= shift_reg_42_im;
    shift_reg_44_re <= shift_reg_43_re;
    shift_reg_44_im <= shift_reg_43_im;
    shift_reg_45_re <= shift_reg_44_re;
    shift_reg_45_im <= shift_reg_44_im;
    shift_reg_46_re <= shift_reg_45_re;
    shift_reg_46_im <= shift_reg_45_im;
    shift_reg_47_re <= shift_reg_46_re;
    shift_reg_47_im <= shift_reg_46_im;
    shift_reg_48_re <= shift_reg_47_re;
    shift_reg_48_im <= shift_reg_47_im;
    shift_reg_49_re <= shift_reg_48_re;
    shift_reg_49_im <= shift_reg_48_im;
    shift_reg_50_re <= shift_reg_49_re;
    shift_reg_50_im <= shift_reg_49_im;
    shift_reg_51_re <= shift_reg_50_re;
    shift_reg_51_im <= shift_reg_50_im;
    shift_reg_52_re <= shift_reg_51_re;
    shift_reg_52_im <= shift_reg_51_im;
    shift_reg_53_re <= shift_reg_52_re;
    shift_reg_53_im <= shift_reg_52_im;
    shift_reg_54_re <= shift_reg_53_re;
    shift_reg_54_im <= shift_reg_53_im;
    shift_reg_55_re <= shift_reg_54_re;
    shift_reg_55_im <= shift_reg_54_im;
    shift_reg_56_re <= shift_reg_55_re;
    shift_reg_56_im <= shift_reg_55_im;
    shift_reg_57_re <= shift_reg_56_re;
    shift_reg_57_im <= shift_reg_56_im;
    shift_reg_58_re <= shift_reg_57_re;
    shift_reg_58_im <= shift_reg_57_im;
    shift_reg_59_re <= shift_reg_58_re;
    shift_reg_59_im <= shift_reg_58_im;
    shift_reg_60_re <= shift_reg_59_re;
    shift_reg_60_im <= shift_reg_59_im;
    shift_reg_61_re <= shift_reg_60_re;
    shift_reg_61_im <= shift_reg_60_im;
    shift_reg_62_re <= shift_reg_61_re;
    shift_reg_62_im <= shift_reg_61_im;
    shift_reg_63_re <= shift_reg_62_re;
    shift_reg_63_im <= shift_reg_62_im;
  end


endmodule

//R2Butterfly replaced by R2Butterfly

//ShiftRegisterNE_5 replaced by ShiftRegisterNE_5

//R2Switch replaced by R2Switch

module ShiftRegisterNE_5 (
  input      [23:0]   input_re,
  input      [23:0]   input_im,
  output     [23:0]   output_re,
  output     [23:0]   output_im,
  input               clk,
  input               reset
);
  reg        [23:0]   shift_reg_0_re;
  reg        [23:0]   shift_reg_0_im;
  reg        [23:0]   shift_reg_1_re;
  reg        [23:0]   shift_reg_1_im;
  reg        [23:0]   shift_reg_2_re;
  reg        [23:0]   shift_reg_2_im;
  reg        [23:0]   shift_reg_3_re;
  reg        [23:0]   shift_reg_3_im;
  reg        [23:0]   shift_reg_4_re;
  reg        [23:0]   shift_reg_4_im;
  reg        [23:0]   shift_reg_5_re;
  reg        [23:0]   shift_reg_5_im;
  reg        [23:0]   shift_reg_6_re;
  reg        [23:0]   shift_reg_6_im;
  reg        [23:0]   shift_reg_7_re;
  reg        [23:0]   shift_reg_7_im;
  reg        [23:0]   shift_reg_8_re;
  reg        [23:0]   shift_reg_8_im;
  reg        [23:0]   shift_reg_9_re;
  reg        [23:0]   shift_reg_9_im;
  reg        [23:0]   shift_reg_10_re;
  reg        [23:0]   shift_reg_10_im;
  reg        [23:0]   shift_reg_11_re;
  reg        [23:0]   shift_reg_11_im;
  reg        [23:0]   shift_reg_12_re;
  reg        [23:0]   shift_reg_12_im;
  reg        [23:0]   shift_reg_13_re;
  reg        [23:0]   shift_reg_13_im;
  reg        [23:0]   shift_reg_14_re;
  reg        [23:0]   shift_reg_14_im;
  reg        [23:0]   shift_reg_15_re;
  reg        [23:0]   shift_reg_15_im;
  reg        [23:0]   shift_reg_16_re;
  reg        [23:0]   shift_reg_16_im;
  reg        [23:0]   shift_reg_17_re;
  reg        [23:0]   shift_reg_17_im;
  reg        [23:0]   shift_reg_18_re;
  reg        [23:0]   shift_reg_18_im;
  reg        [23:0]   shift_reg_19_re;
  reg        [23:0]   shift_reg_19_im;
  reg        [23:0]   shift_reg_20_re;
  reg        [23:0]   shift_reg_20_im;
  reg        [23:0]   shift_reg_21_re;
  reg        [23:0]   shift_reg_21_im;
  reg        [23:0]   shift_reg_22_re;
  reg        [23:0]   shift_reg_22_im;
  reg        [23:0]   shift_reg_23_re;
  reg        [23:0]   shift_reg_23_im;
  reg        [23:0]   shift_reg_24_re;
  reg        [23:0]   shift_reg_24_im;
  reg        [23:0]   shift_reg_25_re;
  reg        [23:0]   shift_reg_25_im;
  reg        [23:0]   shift_reg_26_re;
  reg        [23:0]   shift_reg_26_im;
  reg        [23:0]   shift_reg_27_re;
  reg        [23:0]   shift_reg_27_im;
  reg        [23:0]   shift_reg_28_re;
  reg        [23:0]   shift_reg_28_im;
  reg        [23:0]   shift_reg_29_re;
  reg        [23:0]   shift_reg_29_im;
  reg        [23:0]   shift_reg_30_re;
  reg        [23:0]   shift_reg_30_im;
  reg        [23:0]   shift_reg_31_re;
  reg        [23:0]   shift_reg_31_im;
  reg        [23:0]   shift_reg_32_re;
  reg        [23:0]   shift_reg_32_im;
  reg        [23:0]   shift_reg_33_re;
  reg        [23:0]   shift_reg_33_im;
  reg        [23:0]   shift_reg_34_re;
  reg        [23:0]   shift_reg_34_im;
  reg        [23:0]   shift_reg_35_re;
  reg        [23:0]   shift_reg_35_im;
  reg        [23:0]   shift_reg_36_re;
  reg        [23:0]   shift_reg_36_im;
  reg        [23:0]   shift_reg_37_re;
  reg        [23:0]   shift_reg_37_im;
  reg        [23:0]   shift_reg_38_re;
  reg        [23:0]   shift_reg_38_im;
  reg        [23:0]   shift_reg_39_re;
  reg        [23:0]   shift_reg_39_im;
  reg        [23:0]   shift_reg_40_re;
  reg        [23:0]   shift_reg_40_im;
  reg        [23:0]   shift_reg_41_re;
  reg        [23:0]   shift_reg_41_im;
  reg        [23:0]   shift_reg_42_re;
  reg        [23:0]   shift_reg_42_im;
  reg        [23:0]   shift_reg_43_re;
  reg        [23:0]   shift_reg_43_im;
  reg        [23:0]   shift_reg_44_re;
  reg        [23:0]   shift_reg_44_im;
  reg        [23:0]   shift_reg_45_re;
  reg        [23:0]   shift_reg_45_im;
  reg        [23:0]   shift_reg_46_re;
  reg        [23:0]   shift_reg_46_im;
  reg        [23:0]   shift_reg_47_re;
  reg        [23:0]   shift_reg_47_im;
  reg        [23:0]   shift_reg_48_re;
  reg        [23:0]   shift_reg_48_im;
  reg        [23:0]   shift_reg_49_re;
  reg        [23:0]   shift_reg_49_im;
  reg        [23:0]   shift_reg_50_re;
  reg        [23:0]   shift_reg_50_im;
  reg        [23:0]   shift_reg_51_re;
  reg        [23:0]   shift_reg_51_im;
  reg        [23:0]   shift_reg_52_re;
  reg        [23:0]   shift_reg_52_im;
  reg        [23:0]   shift_reg_53_re;
  reg        [23:0]   shift_reg_53_im;
  reg        [23:0]   shift_reg_54_re;
  reg        [23:0]   shift_reg_54_im;
  reg        [23:0]   shift_reg_55_re;
  reg        [23:0]   shift_reg_55_im;
  reg        [23:0]   shift_reg_56_re;
  reg        [23:0]   shift_reg_56_im;
  reg        [23:0]   shift_reg_57_re;
  reg        [23:0]   shift_reg_57_im;
  reg        [23:0]   shift_reg_58_re;
  reg        [23:0]   shift_reg_58_im;
  reg        [23:0]   shift_reg_59_re;
  reg        [23:0]   shift_reg_59_im;
  reg        [23:0]   shift_reg_60_re;
  reg        [23:0]   shift_reg_60_im;
  reg        [23:0]   shift_reg_61_re;
  reg        [23:0]   shift_reg_61_im;
  reg        [23:0]   shift_reg_62_re;
  reg        [23:0]   shift_reg_62_im;
  reg        [23:0]   shift_reg_63_re;
  reg        [23:0]   shift_reg_63_im;
  reg        [23:0]   shift_reg_64_re;
  reg        [23:0]   shift_reg_64_im;
  reg        [23:0]   shift_reg_65_re;
  reg        [23:0]   shift_reg_65_im;
  reg        [23:0]   shift_reg_66_re;
  reg        [23:0]   shift_reg_66_im;
  reg        [23:0]   shift_reg_67_re;
  reg        [23:0]   shift_reg_67_im;
  reg        [23:0]   shift_reg_68_re;
  reg        [23:0]   shift_reg_68_im;
  reg        [23:0]   shift_reg_69_re;
  reg        [23:0]   shift_reg_69_im;
  reg        [23:0]   shift_reg_70_re;
  reg        [23:0]   shift_reg_70_im;
  reg        [23:0]   shift_reg_71_re;
  reg        [23:0]   shift_reg_71_im;
  reg        [23:0]   shift_reg_72_re;
  reg        [23:0]   shift_reg_72_im;
  reg        [23:0]   shift_reg_73_re;
  reg        [23:0]   shift_reg_73_im;
  reg        [23:0]   shift_reg_74_re;
  reg        [23:0]   shift_reg_74_im;
  reg        [23:0]   shift_reg_75_re;
  reg        [23:0]   shift_reg_75_im;
  reg        [23:0]   shift_reg_76_re;
  reg        [23:0]   shift_reg_76_im;
  reg        [23:0]   shift_reg_77_re;
  reg        [23:0]   shift_reg_77_im;
  reg        [23:0]   shift_reg_78_re;
  reg        [23:0]   shift_reg_78_im;
  reg        [23:0]   shift_reg_79_re;
  reg        [23:0]   shift_reg_79_im;
  reg        [23:0]   shift_reg_80_re;
  reg        [23:0]   shift_reg_80_im;
  reg        [23:0]   shift_reg_81_re;
  reg        [23:0]   shift_reg_81_im;
  reg        [23:0]   shift_reg_82_re;
  reg        [23:0]   shift_reg_82_im;
  reg        [23:0]   shift_reg_83_re;
  reg        [23:0]   shift_reg_83_im;
  reg        [23:0]   shift_reg_84_re;
  reg        [23:0]   shift_reg_84_im;
  reg        [23:0]   shift_reg_85_re;
  reg        [23:0]   shift_reg_85_im;
  reg        [23:0]   shift_reg_86_re;
  reg        [23:0]   shift_reg_86_im;
  reg        [23:0]   shift_reg_87_re;
  reg        [23:0]   shift_reg_87_im;
  reg        [23:0]   shift_reg_88_re;
  reg        [23:0]   shift_reg_88_im;
  reg        [23:0]   shift_reg_89_re;
  reg        [23:0]   shift_reg_89_im;
  reg        [23:0]   shift_reg_90_re;
  reg        [23:0]   shift_reg_90_im;
  reg        [23:0]   shift_reg_91_re;
  reg        [23:0]   shift_reg_91_im;
  reg        [23:0]   shift_reg_92_re;
  reg        [23:0]   shift_reg_92_im;
  reg        [23:0]   shift_reg_93_re;
  reg        [23:0]   shift_reg_93_im;
  reg        [23:0]   shift_reg_94_re;
  reg        [23:0]   shift_reg_94_im;
  reg        [23:0]   shift_reg_95_re;
  reg        [23:0]   shift_reg_95_im;
  reg        [23:0]   shift_reg_96_re;
  reg        [23:0]   shift_reg_96_im;
  reg        [23:0]   shift_reg_97_re;
  reg        [23:0]   shift_reg_97_im;
  reg        [23:0]   shift_reg_98_re;
  reg        [23:0]   shift_reg_98_im;
  reg        [23:0]   shift_reg_99_re;
  reg        [23:0]   shift_reg_99_im;
  reg        [23:0]   shift_reg_100_re;
  reg        [23:0]   shift_reg_100_im;
  reg        [23:0]   shift_reg_101_re;
  reg        [23:0]   shift_reg_101_im;
  reg        [23:0]   shift_reg_102_re;
  reg        [23:0]   shift_reg_102_im;
  reg        [23:0]   shift_reg_103_re;
  reg        [23:0]   shift_reg_103_im;
  reg        [23:0]   shift_reg_104_re;
  reg        [23:0]   shift_reg_104_im;
  reg        [23:0]   shift_reg_105_re;
  reg        [23:0]   shift_reg_105_im;
  reg        [23:0]   shift_reg_106_re;
  reg        [23:0]   shift_reg_106_im;
  reg        [23:0]   shift_reg_107_re;
  reg        [23:0]   shift_reg_107_im;
  reg        [23:0]   shift_reg_108_re;
  reg        [23:0]   shift_reg_108_im;
  reg        [23:0]   shift_reg_109_re;
  reg        [23:0]   shift_reg_109_im;
  reg        [23:0]   shift_reg_110_re;
  reg        [23:0]   shift_reg_110_im;
  reg        [23:0]   shift_reg_111_re;
  reg        [23:0]   shift_reg_111_im;
  reg        [23:0]   shift_reg_112_re;
  reg        [23:0]   shift_reg_112_im;
  reg        [23:0]   shift_reg_113_re;
  reg        [23:0]   shift_reg_113_im;
  reg        [23:0]   shift_reg_114_re;
  reg        [23:0]   shift_reg_114_im;
  reg        [23:0]   shift_reg_115_re;
  reg        [23:0]   shift_reg_115_im;
  reg        [23:0]   shift_reg_116_re;
  reg        [23:0]   shift_reg_116_im;
  reg        [23:0]   shift_reg_117_re;
  reg        [23:0]   shift_reg_117_im;
  reg        [23:0]   shift_reg_118_re;
  reg        [23:0]   shift_reg_118_im;
  reg        [23:0]   shift_reg_119_re;
  reg        [23:0]   shift_reg_119_im;
  reg        [23:0]   shift_reg_120_re;
  reg        [23:0]   shift_reg_120_im;
  reg        [23:0]   shift_reg_121_re;
  reg        [23:0]   shift_reg_121_im;
  reg        [23:0]   shift_reg_122_re;
  reg        [23:0]   shift_reg_122_im;
  reg        [23:0]   shift_reg_123_re;
  reg        [23:0]   shift_reg_123_im;
  reg        [23:0]   shift_reg_124_re;
  reg        [23:0]   shift_reg_124_im;
  reg        [23:0]   shift_reg_125_re;
  reg        [23:0]   shift_reg_125_im;
  reg        [23:0]   shift_reg_126_re;
  reg        [23:0]   shift_reg_126_im;
  reg        [23:0]   shift_reg_127_re;
  reg        [23:0]   shift_reg_127_im;

  assign output_re = shift_reg_127_re;
  assign output_im = shift_reg_127_im;
  always @(posedge clk) begin
    shift_reg_0_re <= input_re;
    shift_reg_0_im <= input_im;
    shift_reg_1_re <= shift_reg_0_re;
    shift_reg_1_im <= shift_reg_0_im;
    shift_reg_2_re <= shift_reg_1_re;
    shift_reg_2_im <= shift_reg_1_im;
    shift_reg_3_re <= shift_reg_2_re;
    shift_reg_3_im <= shift_reg_2_im;
    shift_reg_4_re <= shift_reg_3_re;
    shift_reg_4_im <= shift_reg_3_im;
    shift_reg_5_re <= shift_reg_4_re;
    shift_reg_5_im <= shift_reg_4_im;
    shift_reg_6_re <= shift_reg_5_re;
    shift_reg_6_im <= shift_reg_5_im;
    shift_reg_7_re <= shift_reg_6_re;
    shift_reg_7_im <= shift_reg_6_im;
    shift_reg_8_re <= shift_reg_7_re;
    shift_reg_8_im <= shift_reg_7_im;
    shift_reg_9_re <= shift_reg_8_re;
    shift_reg_9_im <= shift_reg_8_im;
    shift_reg_10_re <= shift_reg_9_re;
    shift_reg_10_im <= shift_reg_9_im;
    shift_reg_11_re <= shift_reg_10_re;
    shift_reg_11_im <= shift_reg_10_im;
    shift_reg_12_re <= shift_reg_11_re;
    shift_reg_12_im <= shift_reg_11_im;
    shift_reg_13_re <= shift_reg_12_re;
    shift_reg_13_im <= shift_reg_12_im;
    shift_reg_14_re <= shift_reg_13_re;
    shift_reg_14_im <= shift_reg_13_im;
    shift_reg_15_re <= shift_reg_14_re;
    shift_reg_15_im <= shift_reg_14_im;
    shift_reg_16_re <= shift_reg_15_re;
    shift_reg_16_im <= shift_reg_15_im;
    shift_reg_17_re <= shift_reg_16_re;
    shift_reg_17_im <= shift_reg_16_im;
    shift_reg_18_re <= shift_reg_17_re;
    shift_reg_18_im <= shift_reg_17_im;
    shift_reg_19_re <= shift_reg_18_re;
    shift_reg_19_im <= shift_reg_18_im;
    shift_reg_20_re <= shift_reg_19_re;
    shift_reg_20_im <= shift_reg_19_im;
    shift_reg_21_re <= shift_reg_20_re;
    shift_reg_21_im <= shift_reg_20_im;
    shift_reg_22_re <= shift_reg_21_re;
    shift_reg_22_im <= shift_reg_21_im;
    shift_reg_23_re <= shift_reg_22_re;
    shift_reg_23_im <= shift_reg_22_im;
    shift_reg_24_re <= shift_reg_23_re;
    shift_reg_24_im <= shift_reg_23_im;
    shift_reg_25_re <= shift_reg_24_re;
    shift_reg_25_im <= shift_reg_24_im;
    shift_reg_26_re <= shift_reg_25_re;
    shift_reg_26_im <= shift_reg_25_im;
    shift_reg_27_re <= shift_reg_26_re;
    shift_reg_27_im <= shift_reg_26_im;
    shift_reg_28_re <= shift_reg_27_re;
    shift_reg_28_im <= shift_reg_27_im;
    shift_reg_29_re <= shift_reg_28_re;
    shift_reg_29_im <= shift_reg_28_im;
    shift_reg_30_re <= shift_reg_29_re;
    shift_reg_30_im <= shift_reg_29_im;
    shift_reg_31_re <= shift_reg_30_re;
    shift_reg_31_im <= shift_reg_30_im;
    shift_reg_32_re <= shift_reg_31_re;
    shift_reg_32_im <= shift_reg_31_im;
    shift_reg_33_re <= shift_reg_32_re;
    shift_reg_33_im <= shift_reg_32_im;
    shift_reg_34_re <= shift_reg_33_re;
    shift_reg_34_im <= shift_reg_33_im;
    shift_reg_35_re <= shift_reg_34_re;
    shift_reg_35_im <= shift_reg_34_im;
    shift_reg_36_re <= shift_reg_35_re;
    shift_reg_36_im <= shift_reg_35_im;
    shift_reg_37_re <= shift_reg_36_re;
    shift_reg_37_im <= shift_reg_36_im;
    shift_reg_38_re <= shift_reg_37_re;
    shift_reg_38_im <= shift_reg_37_im;
    shift_reg_39_re <= shift_reg_38_re;
    shift_reg_39_im <= shift_reg_38_im;
    shift_reg_40_re <= shift_reg_39_re;
    shift_reg_40_im <= shift_reg_39_im;
    shift_reg_41_re <= shift_reg_40_re;
    shift_reg_41_im <= shift_reg_40_im;
    shift_reg_42_re <= shift_reg_41_re;
    shift_reg_42_im <= shift_reg_41_im;
    shift_reg_43_re <= shift_reg_42_re;
    shift_reg_43_im <= shift_reg_42_im;
    shift_reg_44_re <= shift_reg_43_re;
    shift_reg_44_im <= shift_reg_43_im;
    shift_reg_45_re <= shift_reg_44_re;
    shift_reg_45_im <= shift_reg_44_im;
    shift_reg_46_re <= shift_reg_45_re;
    shift_reg_46_im <= shift_reg_45_im;
    shift_reg_47_re <= shift_reg_46_re;
    shift_reg_47_im <= shift_reg_46_im;
    shift_reg_48_re <= shift_reg_47_re;
    shift_reg_48_im <= shift_reg_47_im;
    shift_reg_49_re <= shift_reg_48_re;
    shift_reg_49_im <= shift_reg_48_im;
    shift_reg_50_re <= shift_reg_49_re;
    shift_reg_50_im <= shift_reg_49_im;
    shift_reg_51_re <= shift_reg_50_re;
    shift_reg_51_im <= shift_reg_50_im;
    shift_reg_52_re <= shift_reg_51_re;
    shift_reg_52_im <= shift_reg_51_im;
    shift_reg_53_re <= shift_reg_52_re;
    shift_reg_53_im <= shift_reg_52_im;
    shift_reg_54_re <= shift_reg_53_re;
    shift_reg_54_im <= shift_reg_53_im;
    shift_reg_55_re <= shift_reg_54_re;
    shift_reg_55_im <= shift_reg_54_im;
    shift_reg_56_re <= shift_reg_55_re;
    shift_reg_56_im <= shift_reg_55_im;
    shift_reg_57_re <= shift_reg_56_re;
    shift_reg_57_im <= shift_reg_56_im;
    shift_reg_58_re <= shift_reg_57_re;
    shift_reg_58_im <= shift_reg_57_im;
    shift_reg_59_re <= shift_reg_58_re;
    shift_reg_59_im <= shift_reg_58_im;
    shift_reg_60_re <= shift_reg_59_re;
    shift_reg_60_im <= shift_reg_59_im;
    shift_reg_61_re <= shift_reg_60_re;
    shift_reg_61_im <= shift_reg_60_im;
    shift_reg_62_re <= shift_reg_61_re;
    shift_reg_62_im <= shift_reg_61_im;
    shift_reg_63_re <= shift_reg_62_re;
    shift_reg_63_im <= shift_reg_62_im;
    shift_reg_64_re <= shift_reg_63_re;
    shift_reg_64_im <= shift_reg_63_im;
    shift_reg_65_re <= shift_reg_64_re;
    shift_reg_65_im <= shift_reg_64_im;
    shift_reg_66_re <= shift_reg_65_re;
    shift_reg_66_im <= shift_reg_65_im;
    shift_reg_67_re <= shift_reg_66_re;
    shift_reg_67_im <= shift_reg_66_im;
    shift_reg_68_re <= shift_reg_67_re;
    shift_reg_68_im <= shift_reg_67_im;
    shift_reg_69_re <= shift_reg_68_re;
    shift_reg_69_im <= shift_reg_68_im;
    shift_reg_70_re <= shift_reg_69_re;
    shift_reg_70_im <= shift_reg_69_im;
    shift_reg_71_re <= shift_reg_70_re;
    shift_reg_71_im <= shift_reg_70_im;
    shift_reg_72_re <= shift_reg_71_re;
    shift_reg_72_im <= shift_reg_71_im;
    shift_reg_73_re <= shift_reg_72_re;
    shift_reg_73_im <= shift_reg_72_im;
    shift_reg_74_re <= shift_reg_73_re;
    shift_reg_74_im <= shift_reg_73_im;
    shift_reg_75_re <= shift_reg_74_re;
    shift_reg_75_im <= shift_reg_74_im;
    shift_reg_76_re <= shift_reg_75_re;
    shift_reg_76_im <= shift_reg_75_im;
    shift_reg_77_re <= shift_reg_76_re;
    shift_reg_77_im <= shift_reg_76_im;
    shift_reg_78_re <= shift_reg_77_re;
    shift_reg_78_im <= shift_reg_77_im;
    shift_reg_79_re <= shift_reg_78_re;
    shift_reg_79_im <= shift_reg_78_im;
    shift_reg_80_re <= shift_reg_79_re;
    shift_reg_80_im <= shift_reg_79_im;
    shift_reg_81_re <= shift_reg_80_re;
    shift_reg_81_im <= shift_reg_80_im;
    shift_reg_82_re <= shift_reg_81_re;
    shift_reg_82_im <= shift_reg_81_im;
    shift_reg_83_re <= shift_reg_82_re;
    shift_reg_83_im <= shift_reg_82_im;
    shift_reg_84_re <= shift_reg_83_re;
    shift_reg_84_im <= shift_reg_83_im;
    shift_reg_85_re <= shift_reg_84_re;
    shift_reg_85_im <= shift_reg_84_im;
    shift_reg_86_re <= shift_reg_85_re;
    shift_reg_86_im <= shift_reg_85_im;
    shift_reg_87_re <= shift_reg_86_re;
    shift_reg_87_im <= shift_reg_86_im;
    shift_reg_88_re <= shift_reg_87_re;
    shift_reg_88_im <= shift_reg_87_im;
    shift_reg_89_re <= shift_reg_88_re;
    shift_reg_89_im <= shift_reg_88_im;
    shift_reg_90_re <= shift_reg_89_re;
    shift_reg_90_im <= shift_reg_89_im;
    shift_reg_91_re <= shift_reg_90_re;
    shift_reg_91_im <= shift_reg_90_im;
    shift_reg_92_re <= shift_reg_91_re;
    shift_reg_92_im <= shift_reg_91_im;
    shift_reg_93_re <= shift_reg_92_re;
    shift_reg_93_im <= shift_reg_92_im;
    shift_reg_94_re <= shift_reg_93_re;
    shift_reg_94_im <= shift_reg_93_im;
    shift_reg_95_re <= shift_reg_94_re;
    shift_reg_95_im <= shift_reg_94_im;
    shift_reg_96_re <= shift_reg_95_re;
    shift_reg_96_im <= shift_reg_95_im;
    shift_reg_97_re <= shift_reg_96_re;
    shift_reg_97_im <= shift_reg_96_im;
    shift_reg_98_re <= shift_reg_97_re;
    shift_reg_98_im <= shift_reg_97_im;
    shift_reg_99_re <= shift_reg_98_re;
    shift_reg_99_im <= shift_reg_98_im;
    shift_reg_100_re <= shift_reg_99_re;
    shift_reg_100_im <= shift_reg_99_im;
    shift_reg_101_re <= shift_reg_100_re;
    shift_reg_101_im <= shift_reg_100_im;
    shift_reg_102_re <= shift_reg_101_re;
    shift_reg_102_im <= shift_reg_101_im;
    shift_reg_103_re <= shift_reg_102_re;
    shift_reg_103_im <= shift_reg_102_im;
    shift_reg_104_re <= shift_reg_103_re;
    shift_reg_104_im <= shift_reg_103_im;
    shift_reg_105_re <= shift_reg_104_re;
    shift_reg_105_im <= shift_reg_104_im;
    shift_reg_106_re <= shift_reg_105_re;
    shift_reg_106_im <= shift_reg_105_im;
    shift_reg_107_re <= shift_reg_106_re;
    shift_reg_107_im <= shift_reg_106_im;
    shift_reg_108_re <= shift_reg_107_re;
    shift_reg_108_im <= shift_reg_107_im;
    shift_reg_109_re <= shift_reg_108_re;
    shift_reg_109_im <= shift_reg_108_im;
    shift_reg_110_re <= shift_reg_109_re;
    shift_reg_110_im <= shift_reg_109_im;
    shift_reg_111_re <= shift_reg_110_re;
    shift_reg_111_im <= shift_reg_110_im;
    shift_reg_112_re <= shift_reg_111_re;
    shift_reg_112_im <= shift_reg_111_im;
    shift_reg_113_re <= shift_reg_112_re;
    shift_reg_113_im <= shift_reg_112_im;
    shift_reg_114_re <= shift_reg_113_re;
    shift_reg_114_im <= shift_reg_113_im;
    shift_reg_115_re <= shift_reg_114_re;
    shift_reg_115_im <= shift_reg_114_im;
    shift_reg_116_re <= shift_reg_115_re;
    shift_reg_116_im <= shift_reg_115_im;
    shift_reg_117_re <= shift_reg_116_re;
    shift_reg_117_im <= shift_reg_116_im;
    shift_reg_118_re <= shift_reg_117_re;
    shift_reg_118_im <= shift_reg_117_im;
    shift_reg_119_re <= shift_reg_118_re;
    shift_reg_119_im <= shift_reg_118_im;
    shift_reg_120_re <= shift_reg_119_re;
    shift_reg_120_im <= shift_reg_119_im;
    shift_reg_121_re <= shift_reg_120_re;
    shift_reg_121_im <= shift_reg_120_im;
    shift_reg_122_re <= shift_reg_121_re;
    shift_reg_122_im <= shift_reg_121_im;
    shift_reg_123_re <= shift_reg_122_re;
    shift_reg_123_im <= shift_reg_122_im;
    shift_reg_124_re <= shift_reg_123_re;
    shift_reg_124_im <= shift_reg_123_im;
    shift_reg_125_re <= shift_reg_124_re;
    shift_reg_125_im <= shift_reg_124_im;
    shift_reg_126_re <= shift_reg_125_re;
    shift_reg_126_im <= shift_reg_125_im;
    shift_reg_127_re <= shift_reg_126_re;
    shift_reg_127_im <= shift_reg_126_im;
  end


endmodule

//R2Butterfly replaced by R2Butterfly

//ShiftRegisterNE_3 replaced by ShiftRegisterNE_3

//R2Switch replaced by R2Switch

module ShiftRegisterNE_3 (
  input      [23:0]   input_re,
  input      [23:0]   input_im,
  output     [23:0]   output_re,
  output     [23:0]   output_im,
  input               clk,
  input               reset
);
  reg        [23:0]   shift_reg_0_re;
  reg        [23:0]   shift_reg_0_im;
  reg        [23:0]   shift_reg_1_re;
  reg        [23:0]   shift_reg_1_im;
  reg        [23:0]   shift_reg_2_re;
  reg        [23:0]   shift_reg_2_im;
  reg        [23:0]   shift_reg_3_re;
  reg        [23:0]   shift_reg_3_im;
  reg        [23:0]   shift_reg_4_re;
  reg        [23:0]   shift_reg_4_im;
  reg        [23:0]   shift_reg_5_re;
  reg        [23:0]   shift_reg_5_im;
  reg        [23:0]   shift_reg_6_re;
  reg        [23:0]   shift_reg_6_im;
  reg        [23:0]   shift_reg_7_re;
  reg        [23:0]   shift_reg_7_im;
  reg        [23:0]   shift_reg_8_re;
  reg        [23:0]   shift_reg_8_im;
  reg        [23:0]   shift_reg_9_re;
  reg        [23:0]   shift_reg_9_im;
  reg        [23:0]   shift_reg_10_re;
  reg        [23:0]   shift_reg_10_im;
  reg        [23:0]   shift_reg_11_re;
  reg        [23:0]   shift_reg_11_im;
  reg        [23:0]   shift_reg_12_re;
  reg        [23:0]   shift_reg_12_im;
  reg        [23:0]   shift_reg_13_re;
  reg        [23:0]   shift_reg_13_im;
  reg        [23:0]   shift_reg_14_re;
  reg        [23:0]   shift_reg_14_im;
  reg        [23:0]   shift_reg_15_re;
  reg        [23:0]   shift_reg_15_im;
  reg        [23:0]   shift_reg_16_re;
  reg        [23:0]   shift_reg_16_im;
  reg        [23:0]   shift_reg_17_re;
  reg        [23:0]   shift_reg_17_im;
  reg        [23:0]   shift_reg_18_re;
  reg        [23:0]   shift_reg_18_im;
  reg        [23:0]   shift_reg_19_re;
  reg        [23:0]   shift_reg_19_im;
  reg        [23:0]   shift_reg_20_re;
  reg        [23:0]   shift_reg_20_im;
  reg        [23:0]   shift_reg_21_re;
  reg        [23:0]   shift_reg_21_im;
  reg        [23:0]   shift_reg_22_re;
  reg        [23:0]   shift_reg_22_im;
  reg        [23:0]   shift_reg_23_re;
  reg        [23:0]   shift_reg_23_im;
  reg        [23:0]   shift_reg_24_re;
  reg        [23:0]   shift_reg_24_im;
  reg        [23:0]   shift_reg_25_re;
  reg        [23:0]   shift_reg_25_im;
  reg        [23:0]   shift_reg_26_re;
  reg        [23:0]   shift_reg_26_im;
  reg        [23:0]   shift_reg_27_re;
  reg        [23:0]   shift_reg_27_im;
  reg        [23:0]   shift_reg_28_re;
  reg        [23:0]   shift_reg_28_im;
  reg        [23:0]   shift_reg_29_re;
  reg        [23:0]   shift_reg_29_im;
  reg        [23:0]   shift_reg_30_re;
  reg        [23:0]   shift_reg_30_im;
  reg        [23:0]   shift_reg_31_re;
  reg        [23:0]   shift_reg_31_im;
  reg        [23:0]   shift_reg_32_re;
  reg        [23:0]   shift_reg_32_im;
  reg        [23:0]   shift_reg_33_re;
  reg        [23:0]   shift_reg_33_im;
  reg        [23:0]   shift_reg_34_re;
  reg        [23:0]   shift_reg_34_im;
  reg        [23:0]   shift_reg_35_re;
  reg        [23:0]   shift_reg_35_im;
  reg        [23:0]   shift_reg_36_re;
  reg        [23:0]   shift_reg_36_im;
  reg        [23:0]   shift_reg_37_re;
  reg        [23:0]   shift_reg_37_im;
  reg        [23:0]   shift_reg_38_re;
  reg        [23:0]   shift_reg_38_im;
  reg        [23:0]   shift_reg_39_re;
  reg        [23:0]   shift_reg_39_im;
  reg        [23:0]   shift_reg_40_re;
  reg        [23:0]   shift_reg_40_im;
  reg        [23:0]   shift_reg_41_re;
  reg        [23:0]   shift_reg_41_im;
  reg        [23:0]   shift_reg_42_re;
  reg        [23:0]   shift_reg_42_im;
  reg        [23:0]   shift_reg_43_re;
  reg        [23:0]   shift_reg_43_im;
  reg        [23:0]   shift_reg_44_re;
  reg        [23:0]   shift_reg_44_im;
  reg        [23:0]   shift_reg_45_re;
  reg        [23:0]   shift_reg_45_im;
  reg        [23:0]   shift_reg_46_re;
  reg        [23:0]   shift_reg_46_im;
  reg        [23:0]   shift_reg_47_re;
  reg        [23:0]   shift_reg_47_im;
  reg        [23:0]   shift_reg_48_re;
  reg        [23:0]   shift_reg_48_im;
  reg        [23:0]   shift_reg_49_re;
  reg        [23:0]   shift_reg_49_im;
  reg        [23:0]   shift_reg_50_re;
  reg        [23:0]   shift_reg_50_im;
  reg        [23:0]   shift_reg_51_re;
  reg        [23:0]   shift_reg_51_im;
  reg        [23:0]   shift_reg_52_re;
  reg        [23:0]   shift_reg_52_im;
  reg        [23:0]   shift_reg_53_re;
  reg        [23:0]   shift_reg_53_im;
  reg        [23:0]   shift_reg_54_re;
  reg        [23:0]   shift_reg_54_im;
  reg        [23:0]   shift_reg_55_re;
  reg        [23:0]   shift_reg_55_im;
  reg        [23:0]   shift_reg_56_re;
  reg        [23:0]   shift_reg_56_im;
  reg        [23:0]   shift_reg_57_re;
  reg        [23:0]   shift_reg_57_im;
  reg        [23:0]   shift_reg_58_re;
  reg        [23:0]   shift_reg_58_im;
  reg        [23:0]   shift_reg_59_re;
  reg        [23:0]   shift_reg_59_im;
  reg        [23:0]   shift_reg_60_re;
  reg        [23:0]   shift_reg_60_im;
  reg        [23:0]   shift_reg_61_re;
  reg        [23:0]   shift_reg_61_im;
  reg        [23:0]   shift_reg_62_re;
  reg        [23:0]   shift_reg_62_im;
  reg        [23:0]   shift_reg_63_re;
  reg        [23:0]   shift_reg_63_im;
  reg        [23:0]   shift_reg_64_re;
  reg        [23:0]   shift_reg_64_im;
  reg        [23:0]   shift_reg_65_re;
  reg        [23:0]   shift_reg_65_im;
  reg        [23:0]   shift_reg_66_re;
  reg        [23:0]   shift_reg_66_im;
  reg        [23:0]   shift_reg_67_re;
  reg        [23:0]   shift_reg_67_im;
  reg        [23:0]   shift_reg_68_re;
  reg        [23:0]   shift_reg_68_im;
  reg        [23:0]   shift_reg_69_re;
  reg        [23:0]   shift_reg_69_im;
  reg        [23:0]   shift_reg_70_re;
  reg        [23:0]   shift_reg_70_im;
  reg        [23:0]   shift_reg_71_re;
  reg        [23:0]   shift_reg_71_im;
  reg        [23:0]   shift_reg_72_re;
  reg        [23:0]   shift_reg_72_im;
  reg        [23:0]   shift_reg_73_re;
  reg        [23:0]   shift_reg_73_im;
  reg        [23:0]   shift_reg_74_re;
  reg        [23:0]   shift_reg_74_im;
  reg        [23:0]   shift_reg_75_re;
  reg        [23:0]   shift_reg_75_im;
  reg        [23:0]   shift_reg_76_re;
  reg        [23:0]   shift_reg_76_im;
  reg        [23:0]   shift_reg_77_re;
  reg        [23:0]   shift_reg_77_im;
  reg        [23:0]   shift_reg_78_re;
  reg        [23:0]   shift_reg_78_im;
  reg        [23:0]   shift_reg_79_re;
  reg        [23:0]   shift_reg_79_im;
  reg        [23:0]   shift_reg_80_re;
  reg        [23:0]   shift_reg_80_im;
  reg        [23:0]   shift_reg_81_re;
  reg        [23:0]   shift_reg_81_im;
  reg        [23:0]   shift_reg_82_re;
  reg        [23:0]   shift_reg_82_im;
  reg        [23:0]   shift_reg_83_re;
  reg        [23:0]   shift_reg_83_im;
  reg        [23:0]   shift_reg_84_re;
  reg        [23:0]   shift_reg_84_im;
  reg        [23:0]   shift_reg_85_re;
  reg        [23:0]   shift_reg_85_im;
  reg        [23:0]   shift_reg_86_re;
  reg        [23:0]   shift_reg_86_im;
  reg        [23:0]   shift_reg_87_re;
  reg        [23:0]   shift_reg_87_im;
  reg        [23:0]   shift_reg_88_re;
  reg        [23:0]   shift_reg_88_im;
  reg        [23:0]   shift_reg_89_re;
  reg        [23:0]   shift_reg_89_im;
  reg        [23:0]   shift_reg_90_re;
  reg        [23:0]   shift_reg_90_im;
  reg        [23:0]   shift_reg_91_re;
  reg        [23:0]   shift_reg_91_im;
  reg        [23:0]   shift_reg_92_re;
  reg        [23:0]   shift_reg_92_im;
  reg        [23:0]   shift_reg_93_re;
  reg        [23:0]   shift_reg_93_im;
  reg        [23:0]   shift_reg_94_re;
  reg        [23:0]   shift_reg_94_im;
  reg        [23:0]   shift_reg_95_re;
  reg        [23:0]   shift_reg_95_im;
  reg        [23:0]   shift_reg_96_re;
  reg        [23:0]   shift_reg_96_im;
  reg        [23:0]   shift_reg_97_re;
  reg        [23:0]   shift_reg_97_im;
  reg        [23:0]   shift_reg_98_re;
  reg        [23:0]   shift_reg_98_im;
  reg        [23:0]   shift_reg_99_re;
  reg        [23:0]   shift_reg_99_im;
  reg        [23:0]   shift_reg_100_re;
  reg        [23:0]   shift_reg_100_im;
  reg        [23:0]   shift_reg_101_re;
  reg        [23:0]   shift_reg_101_im;
  reg        [23:0]   shift_reg_102_re;
  reg        [23:0]   shift_reg_102_im;
  reg        [23:0]   shift_reg_103_re;
  reg        [23:0]   shift_reg_103_im;
  reg        [23:0]   shift_reg_104_re;
  reg        [23:0]   shift_reg_104_im;
  reg        [23:0]   shift_reg_105_re;
  reg        [23:0]   shift_reg_105_im;
  reg        [23:0]   shift_reg_106_re;
  reg        [23:0]   shift_reg_106_im;
  reg        [23:0]   shift_reg_107_re;
  reg        [23:0]   shift_reg_107_im;
  reg        [23:0]   shift_reg_108_re;
  reg        [23:0]   shift_reg_108_im;
  reg        [23:0]   shift_reg_109_re;
  reg        [23:0]   shift_reg_109_im;
  reg        [23:0]   shift_reg_110_re;
  reg        [23:0]   shift_reg_110_im;
  reg        [23:0]   shift_reg_111_re;
  reg        [23:0]   shift_reg_111_im;
  reg        [23:0]   shift_reg_112_re;
  reg        [23:0]   shift_reg_112_im;
  reg        [23:0]   shift_reg_113_re;
  reg        [23:0]   shift_reg_113_im;
  reg        [23:0]   shift_reg_114_re;
  reg        [23:0]   shift_reg_114_im;
  reg        [23:0]   shift_reg_115_re;
  reg        [23:0]   shift_reg_115_im;
  reg        [23:0]   shift_reg_116_re;
  reg        [23:0]   shift_reg_116_im;
  reg        [23:0]   shift_reg_117_re;
  reg        [23:0]   shift_reg_117_im;
  reg        [23:0]   shift_reg_118_re;
  reg        [23:0]   shift_reg_118_im;
  reg        [23:0]   shift_reg_119_re;
  reg        [23:0]   shift_reg_119_im;
  reg        [23:0]   shift_reg_120_re;
  reg        [23:0]   shift_reg_120_im;
  reg        [23:0]   shift_reg_121_re;
  reg        [23:0]   shift_reg_121_im;
  reg        [23:0]   shift_reg_122_re;
  reg        [23:0]   shift_reg_122_im;
  reg        [23:0]   shift_reg_123_re;
  reg        [23:0]   shift_reg_123_im;
  reg        [23:0]   shift_reg_124_re;
  reg        [23:0]   shift_reg_124_im;
  reg        [23:0]   shift_reg_125_re;
  reg        [23:0]   shift_reg_125_im;
  reg        [23:0]   shift_reg_126_re;
  reg        [23:0]   shift_reg_126_im;
  reg        [23:0]   shift_reg_127_re;
  reg        [23:0]   shift_reg_127_im;
  reg        [23:0]   shift_reg_128_re;
  reg        [23:0]   shift_reg_128_im;
  reg        [23:0]   shift_reg_129_re;
  reg        [23:0]   shift_reg_129_im;
  reg        [23:0]   shift_reg_130_re;
  reg        [23:0]   shift_reg_130_im;
  reg        [23:0]   shift_reg_131_re;
  reg        [23:0]   shift_reg_131_im;
  reg        [23:0]   shift_reg_132_re;
  reg        [23:0]   shift_reg_132_im;
  reg        [23:0]   shift_reg_133_re;
  reg        [23:0]   shift_reg_133_im;
  reg        [23:0]   shift_reg_134_re;
  reg        [23:0]   shift_reg_134_im;
  reg        [23:0]   shift_reg_135_re;
  reg        [23:0]   shift_reg_135_im;
  reg        [23:0]   shift_reg_136_re;
  reg        [23:0]   shift_reg_136_im;
  reg        [23:0]   shift_reg_137_re;
  reg        [23:0]   shift_reg_137_im;
  reg        [23:0]   shift_reg_138_re;
  reg        [23:0]   shift_reg_138_im;
  reg        [23:0]   shift_reg_139_re;
  reg        [23:0]   shift_reg_139_im;
  reg        [23:0]   shift_reg_140_re;
  reg        [23:0]   shift_reg_140_im;
  reg        [23:0]   shift_reg_141_re;
  reg        [23:0]   shift_reg_141_im;
  reg        [23:0]   shift_reg_142_re;
  reg        [23:0]   shift_reg_142_im;
  reg        [23:0]   shift_reg_143_re;
  reg        [23:0]   shift_reg_143_im;
  reg        [23:0]   shift_reg_144_re;
  reg        [23:0]   shift_reg_144_im;
  reg        [23:0]   shift_reg_145_re;
  reg        [23:0]   shift_reg_145_im;
  reg        [23:0]   shift_reg_146_re;
  reg        [23:0]   shift_reg_146_im;
  reg        [23:0]   shift_reg_147_re;
  reg        [23:0]   shift_reg_147_im;
  reg        [23:0]   shift_reg_148_re;
  reg        [23:0]   shift_reg_148_im;
  reg        [23:0]   shift_reg_149_re;
  reg        [23:0]   shift_reg_149_im;
  reg        [23:0]   shift_reg_150_re;
  reg        [23:0]   shift_reg_150_im;
  reg        [23:0]   shift_reg_151_re;
  reg        [23:0]   shift_reg_151_im;
  reg        [23:0]   shift_reg_152_re;
  reg        [23:0]   shift_reg_152_im;
  reg        [23:0]   shift_reg_153_re;
  reg        [23:0]   shift_reg_153_im;
  reg        [23:0]   shift_reg_154_re;
  reg        [23:0]   shift_reg_154_im;
  reg        [23:0]   shift_reg_155_re;
  reg        [23:0]   shift_reg_155_im;
  reg        [23:0]   shift_reg_156_re;
  reg        [23:0]   shift_reg_156_im;
  reg        [23:0]   shift_reg_157_re;
  reg        [23:0]   shift_reg_157_im;
  reg        [23:0]   shift_reg_158_re;
  reg        [23:0]   shift_reg_158_im;
  reg        [23:0]   shift_reg_159_re;
  reg        [23:0]   shift_reg_159_im;
  reg        [23:0]   shift_reg_160_re;
  reg        [23:0]   shift_reg_160_im;
  reg        [23:0]   shift_reg_161_re;
  reg        [23:0]   shift_reg_161_im;
  reg        [23:0]   shift_reg_162_re;
  reg        [23:0]   shift_reg_162_im;
  reg        [23:0]   shift_reg_163_re;
  reg        [23:0]   shift_reg_163_im;
  reg        [23:0]   shift_reg_164_re;
  reg        [23:0]   shift_reg_164_im;
  reg        [23:0]   shift_reg_165_re;
  reg        [23:0]   shift_reg_165_im;
  reg        [23:0]   shift_reg_166_re;
  reg        [23:0]   shift_reg_166_im;
  reg        [23:0]   shift_reg_167_re;
  reg        [23:0]   shift_reg_167_im;
  reg        [23:0]   shift_reg_168_re;
  reg        [23:0]   shift_reg_168_im;
  reg        [23:0]   shift_reg_169_re;
  reg        [23:0]   shift_reg_169_im;
  reg        [23:0]   shift_reg_170_re;
  reg        [23:0]   shift_reg_170_im;
  reg        [23:0]   shift_reg_171_re;
  reg        [23:0]   shift_reg_171_im;
  reg        [23:0]   shift_reg_172_re;
  reg        [23:0]   shift_reg_172_im;
  reg        [23:0]   shift_reg_173_re;
  reg        [23:0]   shift_reg_173_im;
  reg        [23:0]   shift_reg_174_re;
  reg        [23:0]   shift_reg_174_im;
  reg        [23:0]   shift_reg_175_re;
  reg        [23:0]   shift_reg_175_im;
  reg        [23:0]   shift_reg_176_re;
  reg        [23:0]   shift_reg_176_im;
  reg        [23:0]   shift_reg_177_re;
  reg        [23:0]   shift_reg_177_im;
  reg        [23:0]   shift_reg_178_re;
  reg        [23:0]   shift_reg_178_im;
  reg        [23:0]   shift_reg_179_re;
  reg        [23:0]   shift_reg_179_im;
  reg        [23:0]   shift_reg_180_re;
  reg        [23:0]   shift_reg_180_im;
  reg        [23:0]   shift_reg_181_re;
  reg        [23:0]   shift_reg_181_im;
  reg        [23:0]   shift_reg_182_re;
  reg        [23:0]   shift_reg_182_im;
  reg        [23:0]   shift_reg_183_re;
  reg        [23:0]   shift_reg_183_im;
  reg        [23:0]   shift_reg_184_re;
  reg        [23:0]   shift_reg_184_im;
  reg        [23:0]   shift_reg_185_re;
  reg        [23:0]   shift_reg_185_im;
  reg        [23:0]   shift_reg_186_re;
  reg        [23:0]   shift_reg_186_im;
  reg        [23:0]   shift_reg_187_re;
  reg        [23:0]   shift_reg_187_im;
  reg        [23:0]   shift_reg_188_re;
  reg        [23:0]   shift_reg_188_im;
  reg        [23:0]   shift_reg_189_re;
  reg        [23:0]   shift_reg_189_im;
  reg        [23:0]   shift_reg_190_re;
  reg        [23:0]   shift_reg_190_im;
  reg        [23:0]   shift_reg_191_re;
  reg        [23:0]   shift_reg_191_im;
  reg        [23:0]   shift_reg_192_re;
  reg        [23:0]   shift_reg_192_im;
  reg        [23:0]   shift_reg_193_re;
  reg        [23:0]   shift_reg_193_im;
  reg        [23:0]   shift_reg_194_re;
  reg        [23:0]   shift_reg_194_im;
  reg        [23:0]   shift_reg_195_re;
  reg        [23:0]   shift_reg_195_im;
  reg        [23:0]   shift_reg_196_re;
  reg        [23:0]   shift_reg_196_im;
  reg        [23:0]   shift_reg_197_re;
  reg        [23:0]   shift_reg_197_im;
  reg        [23:0]   shift_reg_198_re;
  reg        [23:0]   shift_reg_198_im;
  reg        [23:0]   shift_reg_199_re;
  reg        [23:0]   shift_reg_199_im;
  reg        [23:0]   shift_reg_200_re;
  reg        [23:0]   shift_reg_200_im;
  reg        [23:0]   shift_reg_201_re;
  reg        [23:0]   shift_reg_201_im;
  reg        [23:0]   shift_reg_202_re;
  reg        [23:0]   shift_reg_202_im;
  reg        [23:0]   shift_reg_203_re;
  reg        [23:0]   shift_reg_203_im;
  reg        [23:0]   shift_reg_204_re;
  reg        [23:0]   shift_reg_204_im;
  reg        [23:0]   shift_reg_205_re;
  reg        [23:0]   shift_reg_205_im;
  reg        [23:0]   shift_reg_206_re;
  reg        [23:0]   shift_reg_206_im;
  reg        [23:0]   shift_reg_207_re;
  reg        [23:0]   shift_reg_207_im;
  reg        [23:0]   shift_reg_208_re;
  reg        [23:0]   shift_reg_208_im;
  reg        [23:0]   shift_reg_209_re;
  reg        [23:0]   shift_reg_209_im;
  reg        [23:0]   shift_reg_210_re;
  reg        [23:0]   shift_reg_210_im;
  reg        [23:0]   shift_reg_211_re;
  reg        [23:0]   shift_reg_211_im;
  reg        [23:0]   shift_reg_212_re;
  reg        [23:0]   shift_reg_212_im;
  reg        [23:0]   shift_reg_213_re;
  reg        [23:0]   shift_reg_213_im;
  reg        [23:0]   shift_reg_214_re;
  reg        [23:0]   shift_reg_214_im;
  reg        [23:0]   shift_reg_215_re;
  reg        [23:0]   shift_reg_215_im;
  reg        [23:0]   shift_reg_216_re;
  reg        [23:0]   shift_reg_216_im;
  reg        [23:0]   shift_reg_217_re;
  reg        [23:0]   shift_reg_217_im;
  reg        [23:0]   shift_reg_218_re;
  reg        [23:0]   shift_reg_218_im;
  reg        [23:0]   shift_reg_219_re;
  reg        [23:0]   shift_reg_219_im;
  reg        [23:0]   shift_reg_220_re;
  reg        [23:0]   shift_reg_220_im;
  reg        [23:0]   shift_reg_221_re;
  reg        [23:0]   shift_reg_221_im;
  reg        [23:0]   shift_reg_222_re;
  reg        [23:0]   shift_reg_222_im;
  reg        [23:0]   shift_reg_223_re;
  reg        [23:0]   shift_reg_223_im;
  reg        [23:0]   shift_reg_224_re;
  reg        [23:0]   shift_reg_224_im;
  reg        [23:0]   shift_reg_225_re;
  reg        [23:0]   shift_reg_225_im;
  reg        [23:0]   shift_reg_226_re;
  reg        [23:0]   shift_reg_226_im;
  reg        [23:0]   shift_reg_227_re;
  reg        [23:0]   shift_reg_227_im;
  reg        [23:0]   shift_reg_228_re;
  reg        [23:0]   shift_reg_228_im;
  reg        [23:0]   shift_reg_229_re;
  reg        [23:0]   shift_reg_229_im;
  reg        [23:0]   shift_reg_230_re;
  reg        [23:0]   shift_reg_230_im;
  reg        [23:0]   shift_reg_231_re;
  reg        [23:0]   shift_reg_231_im;
  reg        [23:0]   shift_reg_232_re;
  reg        [23:0]   shift_reg_232_im;
  reg        [23:0]   shift_reg_233_re;
  reg        [23:0]   shift_reg_233_im;
  reg        [23:0]   shift_reg_234_re;
  reg        [23:0]   shift_reg_234_im;
  reg        [23:0]   shift_reg_235_re;
  reg        [23:0]   shift_reg_235_im;
  reg        [23:0]   shift_reg_236_re;
  reg        [23:0]   shift_reg_236_im;
  reg        [23:0]   shift_reg_237_re;
  reg        [23:0]   shift_reg_237_im;
  reg        [23:0]   shift_reg_238_re;
  reg        [23:0]   shift_reg_238_im;
  reg        [23:0]   shift_reg_239_re;
  reg        [23:0]   shift_reg_239_im;
  reg        [23:0]   shift_reg_240_re;
  reg        [23:0]   shift_reg_240_im;
  reg        [23:0]   shift_reg_241_re;
  reg        [23:0]   shift_reg_241_im;
  reg        [23:0]   shift_reg_242_re;
  reg        [23:0]   shift_reg_242_im;
  reg        [23:0]   shift_reg_243_re;
  reg        [23:0]   shift_reg_243_im;
  reg        [23:0]   shift_reg_244_re;
  reg        [23:0]   shift_reg_244_im;
  reg        [23:0]   shift_reg_245_re;
  reg        [23:0]   shift_reg_245_im;
  reg        [23:0]   shift_reg_246_re;
  reg        [23:0]   shift_reg_246_im;
  reg        [23:0]   shift_reg_247_re;
  reg        [23:0]   shift_reg_247_im;
  reg        [23:0]   shift_reg_248_re;
  reg        [23:0]   shift_reg_248_im;
  reg        [23:0]   shift_reg_249_re;
  reg        [23:0]   shift_reg_249_im;
  reg        [23:0]   shift_reg_250_re;
  reg        [23:0]   shift_reg_250_im;
  reg        [23:0]   shift_reg_251_re;
  reg        [23:0]   shift_reg_251_im;
  reg        [23:0]   shift_reg_252_re;
  reg        [23:0]   shift_reg_252_im;
  reg        [23:0]   shift_reg_253_re;
  reg        [23:0]   shift_reg_253_im;
  reg        [23:0]   shift_reg_254_re;
  reg        [23:0]   shift_reg_254_im;
  reg        [23:0]   shift_reg_255_re;
  reg        [23:0]   shift_reg_255_im;

  assign output_re = shift_reg_255_re;
  assign output_im = shift_reg_255_im;
  always @(posedge clk) begin
    shift_reg_0_re <= input_re;
    shift_reg_0_im <= input_im;
    shift_reg_1_re <= shift_reg_0_re;
    shift_reg_1_im <= shift_reg_0_im;
    shift_reg_2_re <= shift_reg_1_re;
    shift_reg_2_im <= shift_reg_1_im;
    shift_reg_3_re <= shift_reg_2_re;
    shift_reg_3_im <= shift_reg_2_im;
    shift_reg_4_re <= shift_reg_3_re;
    shift_reg_4_im <= shift_reg_3_im;
    shift_reg_5_re <= shift_reg_4_re;
    shift_reg_5_im <= shift_reg_4_im;
    shift_reg_6_re <= shift_reg_5_re;
    shift_reg_6_im <= shift_reg_5_im;
    shift_reg_7_re <= shift_reg_6_re;
    shift_reg_7_im <= shift_reg_6_im;
    shift_reg_8_re <= shift_reg_7_re;
    shift_reg_8_im <= shift_reg_7_im;
    shift_reg_9_re <= shift_reg_8_re;
    shift_reg_9_im <= shift_reg_8_im;
    shift_reg_10_re <= shift_reg_9_re;
    shift_reg_10_im <= shift_reg_9_im;
    shift_reg_11_re <= shift_reg_10_re;
    shift_reg_11_im <= shift_reg_10_im;
    shift_reg_12_re <= shift_reg_11_re;
    shift_reg_12_im <= shift_reg_11_im;
    shift_reg_13_re <= shift_reg_12_re;
    shift_reg_13_im <= shift_reg_12_im;
    shift_reg_14_re <= shift_reg_13_re;
    shift_reg_14_im <= shift_reg_13_im;
    shift_reg_15_re <= shift_reg_14_re;
    shift_reg_15_im <= shift_reg_14_im;
    shift_reg_16_re <= shift_reg_15_re;
    shift_reg_16_im <= shift_reg_15_im;
    shift_reg_17_re <= shift_reg_16_re;
    shift_reg_17_im <= shift_reg_16_im;
    shift_reg_18_re <= shift_reg_17_re;
    shift_reg_18_im <= shift_reg_17_im;
    shift_reg_19_re <= shift_reg_18_re;
    shift_reg_19_im <= shift_reg_18_im;
    shift_reg_20_re <= shift_reg_19_re;
    shift_reg_20_im <= shift_reg_19_im;
    shift_reg_21_re <= shift_reg_20_re;
    shift_reg_21_im <= shift_reg_20_im;
    shift_reg_22_re <= shift_reg_21_re;
    shift_reg_22_im <= shift_reg_21_im;
    shift_reg_23_re <= shift_reg_22_re;
    shift_reg_23_im <= shift_reg_22_im;
    shift_reg_24_re <= shift_reg_23_re;
    shift_reg_24_im <= shift_reg_23_im;
    shift_reg_25_re <= shift_reg_24_re;
    shift_reg_25_im <= shift_reg_24_im;
    shift_reg_26_re <= shift_reg_25_re;
    shift_reg_26_im <= shift_reg_25_im;
    shift_reg_27_re <= shift_reg_26_re;
    shift_reg_27_im <= shift_reg_26_im;
    shift_reg_28_re <= shift_reg_27_re;
    shift_reg_28_im <= shift_reg_27_im;
    shift_reg_29_re <= shift_reg_28_re;
    shift_reg_29_im <= shift_reg_28_im;
    shift_reg_30_re <= shift_reg_29_re;
    shift_reg_30_im <= shift_reg_29_im;
    shift_reg_31_re <= shift_reg_30_re;
    shift_reg_31_im <= shift_reg_30_im;
    shift_reg_32_re <= shift_reg_31_re;
    shift_reg_32_im <= shift_reg_31_im;
    shift_reg_33_re <= shift_reg_32_re;
    shift_reg_33_im <= shift_reg_32_im;
    shift_reg_34_re <= shift_reg_33_re;
    shift_reg_34_im <= shift_reg_33_im;
    shift_reg_35_re <= shift_reg_34_re;
    shift_reg_35_im <= shift_reg_34_im;
    shift_reg_36_re <= shift_reg_35_re;
    shift_reg_36_im <= shift_reg_35_im;
    shift_reg_37_re <= shift_reg_36_re;
    shift_reg_37_im <= shift_reg_36_im;
    shift_reg_38_re <= shift_reg_37_re;
    shift_reg_38_im <= shift_reg_37_im;
    shift_reg_39_re <= shift_reg_38_re;
    shift_reg_39_im <= shift_reg_38_im;
    shift_reg_40_re <= shift_reg_39_re;
    shift_reg_40_im <= shift_reg_39_im;
    shift_reg_41_re <= shift_reg_40_re;
    shift_reg_41_im <= shift_reg_40_im;
    shift_reg_42_re <= shift_reg_41_re;
    shift_reg_42_im <= shift_reg_41_im;
    shift_reg_43_re <= shift_reg_42_re;
    shift_reg_43_im <= shift_reg_42_im;
    shift_reg_44_re <= shift_reg_43_re;
    shift_reg_44_im <= shift_reg_43_im;
    shift_reg_45_re <= shift_reg_44_re;
    shift_reg_45_im <= shift_reg_44_im;
    shift_reg_46_re <= shift_reg_45_re;
    shift_reg_46_im <= shift_reg_45_im;
    shift_reg_47_re <= shift_reg_46_re;
    shift_reg_47_im <= shift_reg_46_im;
    shift_reg_48_re <= shift_reg_47_re;
    shift_reg_48_im <= shift_reg_47_im;
    shift_reg_49_re <= shift_reg_48_re;
    shift_reg_49_im <= shift_reg_48_im;
    shift_reg_50_re <= shift_reg_49_re;
    shift_reg_50_im <= shift_reg_49_im;
    shift_reg_51_re <= shift_reg_50_re;
    shift_reg_51_im <= shift_reg_50_im;
    shift_reg_52_re <= shift_reg_51_re;
    shift_reg_52_im <= shift_reg_51_im;
    shift_reg_53_re <= shift_reg_52_re;
    shift_reg_53_im <= shift_reg_52_im;
    shift_reg_54_re <= shift_reg_53_re;
    shift_reg_54_im <= shift_reg_53_im;
    shift_reg_55_re <= shift_reg_54_re;
    shift_reg_55_im <= shift_reg_54_im;
    shift_reg_56_re <= shift_reg_55_re;
    shift_reg_56_im <= shift_reg_55_im;
    shift_reg_57_re <= shift_reg_56_re;
    shift_reg_57_im <= shift_reg_56_im;
    shift_reg_58_re <= shift_reg_57_re;
    shift_reg_58_im <= shift_reg_57_im;
    shift_reg_59_re <= shift_reg_58_re;
    shift_reg_59_im <= shift_reg_58_im;
    shift_reg_60_re <= shift_reg_59_re;
    shift_reg_60_im <= shift_reg_59_im;
    shift_reg_61_re <= shift_reg_60_re;
    shift_reg_61_im <= shift_reg_60_im;
    shift_reg_62_re <= shift_reg_61_re;
    shift_reg_62_im <= shift_reg_61_im;
    shift_reg_63_re <= shift_reg_62_re;
    shift_reg_63_im <= shift_reg_62_im;
    shift_reg_64_re <= shift_reg_63_re;
    shift_reg_64_im <= shift_reg_63_im;
    shift_reg_65_re <= shift_reg_64_re;
    shift_reg_65_im <= shift_reg_64_im;
    shift_reg_66_re <= shift_reg_65_re;
    shift_reg_66_im <= shift_reg_65_im;
    shift_reg_67_re <= shift_reg_66_re;
    shift_reg_67_im <= shift_reg_66_im;
    shift_reg_68_re <= shift_reg_67_re;
    shift_reg_68_im <= shift_reg_67_im;
    shift_reg_69_re <= shift_reg_68_re;
    shift_reg_69_im <= shift_reg_68_im;
    shift_reg_70_re <= shift_reg_69_re;
    shift_reg_70_im <= shift_reg_69_im;
    shift_reg_71_re <= shift_reg_70_re;
    shift_reg_71_im <= shift_reg_70_im;
    shift_reg_72_re <= shift_reg_71_re;
    shift_reg_72_im <= shift_reg_71_im;
    shift_reg_73_re <= shift_reg_72_re;
    shift_reg_73_im <= shift_reg_72_im;
    shift_reg_74_re <= shift_reg_73_re;
    shift_reg_74_im <= shift_reg_73_im;
    shift_reg_75_re <= shift_reg_74_re;
    shift_reg_75_im <= shift_reg_74_im;
    shift_reg_76_re <= shift_reg_75_re;
    shift_reg_76_im <= shift_reg_75_im;
    shift_reg_77_re <= shift_reg_76_re;
    shift_reg_77_im <= shift_reg_76_im;
    shift_reg_78_re <= shift_reg_77_re;
    shift_reg_78_im <= shift_reg_77_im;
    shift_reg_79_re <= shift_reg_78_re;
    shift_reg_79_im <= shift_reg_78_im;
    shift_reg_80_re <= shift_reg_79_re;
    shift_reg_80_im <= shift_reg_79_im;
    shift_reg_81_re <= shift_reg_80_re;
    shift_reg_81_im <= shift_reg_80_im;
    shift_reg_82_re <= shift_reg_81_re;
    shift_reg_82_im <= shift_reg_81_im;
    shift_reg_83_re <= shift_reg_82_re;
    shift_reg_83_im <= shift_reg_82_im;
    shift_reg_84_re <= shift_reg_83_re;
    shift_reg_84_im <= shift_reg_83_im;
    shift_reg_85_re <= shift_reg_84_re;
    shift_reg_85_im <= shift_reg_84_im;
    shift_reg_86_re <= shift_reg_85_re;
    shift_reg_86_im <= shift_reg_85_im;
    shift_reg_87_re <= shift_reg_86_re;
    shift_reg_87_im <= shift_reg_86_im;
    shift_reg_88_re <= shift_reg_87_re;
    shift_reg_88_im <= shift_reg_87_im;
    shift_reg_89_re <= shift_reg_88_re;
    shift_reg_89_im <= shift_reg_88_im;
    shift_reg_90_re <= shift_reg_89_re;
    shift_reg_90_im <= shift_reg_89_im;
    shift_reg_91_re <= shift_reg_90_re;
    shift_reg_91_im <= shift_reg_90_im;
    shift_reg_92_re <= shift_reg_91_re;
    shift_reg_92_im <= shift_reg_91_im;
    shift_reg_93_re <= shift_reg_92_re;
    shift_reg_93_im <= shift_reg_92_im;
    shift_reg_94_re <= shift_reg_93_re;
    shift_reg_94_im <= shift_reg_93_im;
    shift_reg_95_re <= shift_reg_94_re;
    shift_reg_95_im <= shift_reg_94_im;
    shift_reg_96_re <= shift_reg_95_re;
    shift_reg_96_im <= shift_reg_95_im;
    shift_reg_97_re <= shift_reg_96_re;
    shift_reg_97_im <= shift_reg_96_im;
    shift_reg_98_re <= shift_reg_97_re;
    shift_reg_98_im <= shift_reg_97_im;
    shift_reg_99_re <= shift_reg_98_re;
    shift_reg_99_im <= shift_reg_98_im;
    shift_reg_100_re <= shift_reg_99_re;
    shift_reg_100_im <= shift_reg_99_im;
    shift_reg_101_re <= shift_reg_100_re;
    shift_reg_101_im <= shift_reg_100_im;
    shift_reg_102_re <= shift_reg_101_re;
    shift_reg_102_im <= shift_reg_101_im;
    shift_reg_103_re <= shift_reg_102_re;
    shift_reg_103_im <= shift_reg_102_im;
    shift_reg_104_re <= shift_reg_103_re;
    shift_reg_104_im <= shift_reg_103_im;
    shift_reg_105_re <= shift_reg_104_re;
    shift_reg_105_im <= shift_reg_104_im;
    shift_reg_106_re <= shift_reg_105_re;
    shift_reg_106_im <= shift_reg_105_im;
    shift_reg_107_re <= shift_reg_106_re;
    shift_reg_107_im <= shift_reg_106_im;
    shift_reg_108_re <= shift_reg_107_re;
    shift_reg_108_im <= shift_reg_107_im;
    shift_reg_109_re <= shift_reg_108_re;
    shift_reg_109_im <= shift_reg_108_im;
    shift_reg_110_re <= shift_reg_109_re;
    shift_reg_110_im <= shift_reg_109_im;
    shift_reg_111_re <= shift_reg_110_re;
    shift_reg_111_im <= shift_reg_110_im;
    shift_reg_112_re <= shift_reg_111_re;
    shift_reg_112_im <= shift_reg_111_im;
    shift_reg_113_re <= shift_reg_112_re;
    shift_reg_113_im <= shift_reg_112_im;
    shift_reg_114_re <= shift_reg_113_re;
    shift_reg_114_im <= shift_reg_113_im;
    shift_reg_115_re <= shift_reg_114_re;
    shift_reg_115_im <= shift_reg_114_im;
    shift_reg_116_re <= shift_reg_115_re;
    shift_reg_116_im <= shift_reg_115_im;
    shift_reg_117_re <= shift_reg_116_re;
    shift_reg_117_im <= shift_reg_116_im;
    shift_reg_118_re <= shift_reg_117_re;
    shift_reg_118_im <= shift_reg_117_im;
    shift_reg_119_re <= shift_reg_118_re;
    shift_reg_119_im <= shift_reg_118_im;
    shift_reg_120_re <= shift_reg_119_re;
    shift_reg_120_im <= shift_reg_119_im;
    shift_reg_121_re <= shift_reg_120_re;
    shift_reg_121_im <= shift_reg_120_im;
    shift_reg_122_re <= shift_reg_121_re;
    shift_reg_122_im <= shift_reg_121_im;
    shift_reg_123_re <= shift_reg_122_re;
    shift_reg_123_im <= shift_reg_122_im;
    shift_reg_124_re <= shift_reg_123_re;
    shift_reg_124_im <= shift_reg_123_im;
    shift_reg_125_re <= shift_reg_124_re;
    shift_reg_125_im <= shift_reg_124_im;
    shift_reg_126_re <= shift_reg_125_re;
    shift_reg_126_im <= shift_reg_125_im;
    shift_reg_127_re <= shift_reg_126_re;
    shift_reg_127_im <= shift_reg_126_im;
    shift_reg_128_re <= shift_reg_127_re;
    shift_reg_128_im <= shift_reg_127_im;
    shift_reg_129_re <= shift_reg_128_re;
    shift_reg_129_im <= shift_reg_128_im;
    shift_reg_130_re <= shift_reg_129_re;
    shift_reg_130_im <= shift_reg_129_im;
    shift_reg_131_re <= shift_reg_130_re;
    shift_reg_131_im <= shift_reg_130_im;
    shift_reg_132_re <= shift_reg_131_re;
    shift_reg_132_im <= shift_reg_131_im;
    shift_reg_133_re <= shift_reg_132_re;
    shift_reg_133_im <= shift_reg_132_im;
    shift_reg_134_re <= shift_reg_133_re;
    shift_reg_134_im <= shift_reg_133_im;
    shift_reg_135_re <= shift_reg_134_re;
    shift_reg_135_im <= shift_reg_134_im;
    shift_reg_136_re <= shift_reg_135_re;
    shift_reg_136_im <= shift_reg_135_im;
    shift_reg_137_re <= shift_reg_136_re;
    shift_reg_137_im <= shift_reg_136_im;
    shift_reg_138_re <= shift_reg_137_re;
    shift_reg_138_im <= shift_reg_137_im;
    shift_reg_139_re <= shift_reg_138_re;
    shift_reg_139_im <= shift_reg_138_im;
    shift_reg_140_re <= shift_reg_139_re;
    shift_reg_140_im <= shift_reg_139_im;
    shift_reg_141_re <= shift_reg_140_re;
    shift_reg_141_im <= shift_reg_140_im;
    shift_reg_142_re <= shift_reg_141_re;
    shift_reg_142_im <= shift_reg_141_im;
    shift_reg_143_re <= shift_reg_142_re;
    shift_reg_143_im <= shift_reg_142_im;
    shift_reg_144_re <= shift_reg_143_re;
    shift_reg_144_im <= shift_reg_143_im;
    shift_reg_145_re <= shift_reg_144_re;
    shift_reg_145_im <= shift_reg_144_im;
    shift_reg_146_re <= shift_reg_145_re;
    shift_reg_146_im <= shift_reg_145_im;
    shift_reg_147_re <= shift_reg_146_re;
    shift_reg_147_im <= shift_reg_146_im;
    shift_reg_148_re <= shift_reg_147_re;
    shift_reg_148_im <= shift_reg_147_im;
    shift_reg_149_re <= shift_reg_148_re;
    shift_reg_149_im <= shift_reg_148_im;
    shift_reg_150_re <= shift_reg_149_re;
    shift_reg_150_im <= shift_reg_149_im;
    shift_reg_151_re <= shift_reg_150_re;
    shift_reg_151_im <= shift_reg_150_im;
    shift_reg_152_re <= shift_reg_151_re;
    shift_reg_152_im <= shift_reg_151_im;
    shift_reg_153_re <= shift_reg_152_re;
    shift_reg_153_im <= shift_reg_152_im;
    shift_reg_154_re <= shift_reg_153_re;
    shift_reg_154_im <= shift_reg_153_im;
    shift_reg_155_re <= shift_reg_154_re;
    shift_reg_155_im <= shift_reg_154_im;
    shift_reg_156_re <= shift_reg_155_re;
    shift_reg_156_im <= shift_reg_155_im;
    shift_reg_157_re <= shift_reg_156_re;
    shift_reg_157_im <= shift_reg_156_im;
    shift_reg_158_re <= shift_reg_157_re;
    shift_reg_158_im <= shift_reg_157_im;
    shift_reg_159_re <= shift_reg_158_re;
    shift_reg_159_im <= shift_reg_158_im;
    shift_reg_160_re <= shift_reg_159_re;
    shift_reg_160_im <= shift_reg_159_im;
    shift_reg_161_re <= shift_reg_160_re;
    shift_reg_161_im <= shift_reg_160_im;
    shift_reg_162_re <= shift_reg_161_re;
    shift_reg_162_im <= shift_reg_161_im;
    shift_reg_163_re <= shift_reg_162_re;
    shift_reg_163_im <= shift_reg_162_im;
    shift_reg_164_re <= shift_reg_163_re;
    shift_reg_164_im <= shift_reg_163_im;
    shift_reg_165_re <= shift_reg_164_re;
    shift_reg_165_im <= shift_reg_164_im;
    shift_reg_166_re <= shift_reg_165_re;
    shift_reg_166_im <= shift_reg_165_im;
    shift_reg_167_re <= shift_reg_166_re;
    shift_reg_167_im <= shift_reg_166_im;
    shift_reg_168_re <= shift_reg_167_re;
    shift_reg_168_im <= shift_reg_167_im;
    shift_reg_169_re <= shift_reg_168_re;
    shift_reg_169_im <= shift_reg_168_im;
    shift_reg_170_re <= shift_reg_169_re;
    shift_reg_170_im <= shift_reg_169_im;
    shift_reg_171_re <= shift_reg_170_re;
    shift_reg_171_im <= shift_reg_170_im;
    shift_reg_172_re <= shift_reg_171_re;
    shift_reg_172_im <= shift_reg_171_im;
    shift_reg_173_re <= shift_reg_172_re;
    shift_reg_173_im <= shift_reg_172_im;
    shift_reg_174_re <= shift_reg_173_re;
    shift_reg_174_im <= shift_reg_173_im;
    shift_reg_175_re <= shift_reg_174_re;
    shift_reg_175_im <= shift_reg_174_im;
    shift_reg_176_re <= shift_reg_175_re;
    shift_reg_176_im <= shift_reg_175_im;
    shift_reg_177_re <= shift_reg_176_re;
    shift_reg_177_im <= shift_reg_176_im;
    shift_reg_178_re <= shift_reg_177_re;
    shift_reg_178_im <= shift_reg_177_im;
    shift_reg_179_re <= shift_reg_178_re;
    shift_reg_179_im <= shift_reg_178_im;
    shift_reg_180_re <= shift_reg_179_re;
    shift_reg_180_im <= shift_reg_179_im;
    shift_reg_181_re <= shift_reg_180_re;
    shift_reg_181_im <= shift_reg_180_im;
    shift_reg_182_re <= shift_reg_181_re;
    shift_reg_182_im <= shift_reg_181_im;
    shift_reg_183_re <= shift_reg_182_re;
    shift_reg_183_im <= shift_reg_182_im;
    shift_reg_184_re <= shift_reg_183_re;
    shift_reg_184_im <= shift_reg_183_im;
    shift_reg_185_re <= shift_reg_184_re;
    shift_reg_185_im <= shift_reg_184_im;
    shift_reg_186_re <= shift_reg_185_re;
    shift_reg_186_im <= shift_reg_185_im;
    shift_reg_187_re <= shift_reg_186_re;
    shift_reg_187_im <= shift_reg_186_im;
    shift_reg_188_re <= shift_reg_187_re;
    shift_reg_188_im <= shift_reg_187_im;
    shift_reg_189_re <= shift_reg_188_re;
    shift_reg_189_im <= shift_reg_188_im;
    shift_reg_190_re <= shift_reg_189_re;
    shift_reg_190_im <= shift_reg_189_im;
    shift_reg_191_re <= shift_reg_190_re;
    shift_reg_191_im <= shift_reg_190_im;
    shift_reg_192_re <= shift_reg_191_re;
    shift_reg_192_im <= shift_reg_191_im;
    shift_reg_193_re <= shift_reg_192_re;
    shift_reg_193_im <= shift_reg_192_im;
    shift_reg_194_re <= shift_reg_193_re;
    shift_reg_194_im <= shift_reg_193_im;
    shift_reg_195_re <= shift_reg_194_re;
    shift_reg_195_im <= shift_reg_194_im;
    shift_reg_196_re <= shift_reg_195_re;
    shift_reg_196_im <= shift_reg_195_im;
    shift_reg_197_re <= shift_reg_196_re;
    shift_reg_197_im <= shift_reg_196_im;
    shift_reg_198_re <= shift_reg_197_re;
    shift_reg_198_im <= shift_reg_197_im;
    shift_reg_199_re <= shift_reg_198_re;
    shift_reg_199_im <= shift_reg_198_im;
    shift_reg_200_re <= shift_reg_199_re;
    shift_reg_200_im <= shift_reg_199_im;
    shift_reg_201_re <= shift_reg_200_re;
    shift_reg_201_im <= shift_reg_200_im;
    shift_reg_202_re <= shift_reg_201_re;
    shift_reg_202_im <= shift_reg_201_im;
    shift_reg_203_re <= shift_reg_202_re;
    shift_reg_203_im <= shift_reg_202_im;
    shift_reg_204_re <= shift_reg_203_re;
    shift_reg_204_im <= shift_reg_203_im;
    shift_reg_205_re <= shift_reg_204_re;
    shift_reg_205_im <= shift_reg_204_im;
    shift_reg_206_re <= shift_reg_205_re;
    shift_reg_206_im <= shift_reg_205_im;
    shift_reg_207_re <= shift_reg_206_re;
    shift_reg_207_im <= shift_reg_206_im;
    shift_reg_208_re <= shift_reg_207_re;
    shift_reg_208_im <= shift_reg_207_im;
    shift_reg_209_re <= shift_reg_208_re;
    shift_reg_209_im <= shift_reg_208_im;
    shift_reg_210_re <= shift_reg_209_re;
    shift_reg_210_im <= shift_reg_209_im;
    shift_reg_211_re <= shift_reg_210_re;
    shift_reg_211_im <= shift_reg_210_im;
    shift_reg_212_re <= shift_reg_211_re;
    shift_reg_212_im <= shift_reg_211_im;
    shift_reg_213_re <= shift_reg_212_re;
    shift_reg_213_im <= shift_reg_212_im;
    shift_reg_214_re <= shift_reg_213_re;
    shift_reg_214_im <= shift_reg_213_im;
    shift_reg_215_re <= shift_reg_214_re;
    shift_reg_215_im <= shift_reg_214_im;
    shift_reg_216_re <= shift_reg_215_re;
    shift_reg_216_im <= shift_reg_215_im;
    shift_reg_217_re <= shift_reg_216_re;
    shift_reg_217_im <= shift_reg_216_im;
    shift_reg_218_re <= shift_reg_217_re;
    shift_reg_218_im <= shift_reg_217_im;
    shift_reg_219_re <= shift_reg_218_re;
    shift_reg_219_im <= shift_reg_218_im;
    shift_reg_220_re <= shift_reg_219_re;
    shift_reg_220_im <= shift_reg_219_im;
    shift_reg_221_re <= shift_reg_220_re;
    shift_reg_221_im <= shift_reg_220_im;
    shift_reg_222_re <= shift_reg_221_re;
    shift_reg_222_im <= shift_reg_221_im;
    shift_reg_223_re <= shift_reg_222_re;
    shift_reg_223_im <= shift_reg_222_im;
    shift_reg_224_re <= shift_reg_223_re;
    shift_reg_224_im <= shift_reg_223_im;
    shift_reg_225_re <= shift_reg_224_re;
    shift_reg_225_im <= shift_reg_224_im;
    shift_reg_226_re <= shift_reg_225_re;
    shift_reg_226_im <= shift_reg_225_im;
    shift_reg_227_re <= shift_reg_226_re;
    shift_reg_227_im <= shift_reg_226_im;
    shift_reg_228_re <= shift_reg_227_re;
    shift_reg_228_im <= shift_reg_227_im;
    shift_reg_229_re <= shift_reg_228_re;
    shift_reg_229_im <= shift_reg_228_im;
    shift_reg_230_re <= shift_reg_229_re;
    shift_reg_230_im <= shift_reg_229_im;
    shift_reg_231_re <= shift_reg_230_re;
    shift_reg_231_im <= shift_reg_230_im;
    shift_reg_232_re <= shift_reg_231_re;
    shift_reg_232_im <= shift_reg_231_im;
    shift_reg_233_re <= shift_reg_232_re;
    shift_reg_233_im <= shift_reg_232_im;
    shift_reg_234_re <= shift_reg_233_re;
    shift_reg_234_im <= shift_reg_233_im;
    shift_reg_235_re <= shift_reg_234_re;
    shift_reg_235_im <= shift_reg_234_im;
    shift_reg_236_re <= shift_reg_235_re;
    shift_reg_236_im <= shift_reg_235_im;
    shift_reg_237_re <= shift_reg_236_re;
    shift_reg_237_im <= shift_reg_236_im;
    shift_reg_238_re <= shift_reg_237_re;
    shift_reg_238_im <= shift_reg_237_im;
    shift_reg_239_re <= shift_reg_238_re;
    shift_reg_239_im <= shift_reg_238_im;
    shift_reg_240_re <= shift_reg_239_re;
    shift_reg_240_im <= shift_reg_239_im;
    shift_reg_241_re <= shift_reg_240_re;
    shift_reg_241_im <= shift_reg_240_im;
    shift_reg_242_re <= shift_reg_241_re;
    shift_reg_242_im <= shift_reg_241_im;
    shift_reg_243_re <= shift_reg_242_re;
    shift_reg_243_im <= shift_reg_242_im;
    shift_reg_244_re <= shift_reg_243_re;
    shift_reg_244_im <= shift_reg_243_im;
    shift_reg_245_re <= shift_reg_244_re;
    shift_reg_245_im <= shift_reg_244_im;
    shift_reg_246_re <= shift_reg_245_re;
    shift_reg_246_im <= shift_reg_245_im;
    shift_reg_247_re <= shift_reg_246_re;
    shift_reg_247_im <= shift_reg_246_im;
    shift_reg_248_re <= shift_reg_247_re;
    shift_reg_248_im <= shift_reg_247_im;
    shift_reg_249_re <= shift_reg_248_re;
    shift_reg_249_im <= shift_reg_248_im;
    shift_reg_250_re <= shift_reg_249_re;
    shift_reg_250_im <= shift_reg_249_im;
    shift_reg_251_re <= shift_reg_250_re;
    shift_reg_251_im <= shift_reg_250_im;
    shift_reg_252_re <= shift_reg_251_re;
    shift_reg_252_im <= shift_reg_251_im;
    shift_reg_253_re <= shift_reg_252_re;
    shift_reg_253_im <= shift_reg_252_im;
    shift_reg_254_re <= shift_reg_253_re;
    shift_reg_254_im <= shift_reg_253_im;
    shift_reg_255_re <= shift_reg_254_re;
    shift_reg_255_im <= shift_reg_254_im;
  end


endmodule

//R2Butterfly replaced by R2Butterfly

//ShiftRegisterNE_1 replaced by ShiftRegisterNE_1

module R2Switch (
  input      [23:0]   in1_re,
  input      [23:0]   in1_im,
  input      [23:0]   in2_re,
  input      [23:0]   in2_im,
  input               sel,
  output     [23:0]   out1_re,
  output     [23:0]   out1_im,
  output     [23:0]   out2_re,
  output     [23:0]   out2_im
);

  assign out1_re = (sel ? in2_re : in1_re);
  assign out1_im = (sel ? in2_im : in1_im);
  assign out2_re = (sel ? in1_re : in2_re);
  assign out2_im = (sel ? in1_im : in2_im);

endmodule

module ShiftRegisterNE_1 (
  input      [23:0]   input_re,
  input      [23:0]   input_im,
  output     [23:0]   output_re,
  output     [23:0]   output_im,
  input               clk,
  input               reset
);
  reg        [23:0]   shift_reg_0_re;
  reg        [23:0]   shift_reg_0_im;
  reg        [23:0]   shift_reg_1_re;
  reg        [23:0]   shift_reg_1_im;
  reg        [23:0]   shift_reg_2_re;
  reg        [23:0]   shift_reg_2_im;
  reg        [23:0]   shift_reg_3_re;
  reg        [23:0]   shift_reg_3_im;
  reg        [23:0]   shift_reg_4_re;
  reg        [23:0]   shift_reg_4_im;
  reg        [23:0]   shift_reg_5_re;
  reg        [23:0]   shift_reg_5_im;
  reg        [23:0]   shift_reg_6_re;
  reg        [23:0]   shift_reg_6_im;
  reg        [23:0]   shift_reg_7_re;
  reg        [23:0]   shift_reg_7_im;
  reg        [23:0]   shift_reg_8_re;
  reg        [23:0]   shift_reg_8_im;
  reg        [23:0]   shift_reg_9_re;
  reg        [23:0]   shift_reg_9_im;
  reg        [23:0]   shift_reg_10_re;
  reg        [23:0]   shift_reg_10_im;
  reg        [23:0]   shift_reg_11_re;
  reg        [23:0]   shift_reg_11_im;
  reg        [23:0]   shift_reg_12_re;
  reg        [23:0]   shift_reg_12_im;
  reg        [23:0]   shift_reg_13_re;
  reg        [23:0]   shift_reg_13_im;
  reg        [23:0]   shift_reg_14_re;
  reg        [23:0]   shift_reg_14_im;
  reg        [23:0]   shift_reg_15_re;
  reg        [23:0]   shift_reg_15_im;
  reg        [23:0]   shift_reg_16_re;
  reg        [23:0]   shift_reg_16_im;
  reg        [23:0]   shift_reg_17_re;
  reg        [23:0]   shift_reg_17_im;
  reg        [23:0]   shift_reg_18_re;
  reg        [23:0]   shift_reg_18_im;
  reg        [23:0]   shift_reg_19_re;
  reg        [23:0]   shift_reg_19_im;
  reg        [23:0]   shift_reg_20_re;
  reg        [23:0]   shift_reg_20_im;
  reg        [23:0]   shift_reg_21_re;
  reg        [23:0]   shift_reg_21_im;
  reg        [23:0]   shift_reg_22_re;
  reg        [23:0]   shift_reg_22_im;
  reg        [23:0]   shift_reg_23_re;
  reg        [23:0]   shift_reg_23_im;
  reg        [23:0]   shift_reg_24_re;
  reg        [23:0]   shift_reg_24_im;
  reg        [23:0]   shift_reg_25_re;
  reg        [23:0]   shift_reg_25_im;
  reg        [23:0]   shift_reg_26_re;
  reg        [23:0]   shift_reg_26_im;
  reg        [23:0]   shift_reg_27_re;
  reg        [23:0]   shift_reg_27_im;
  reg        [23:0]   shift_reg_28_re;
  reg        [23:0]   shift_reg_28_im;
  reg        [23:0]   shift_reg_29_re;
  reg        [23:0]   shift_reg_29_im;
  reg        [23:0]   shift_reg_30_re;
  reg        [23:0]   shift_reg_30_im;
  reg        [23:0]   shift_reg_31_re;
  reg        [23:0]   shift_reg_31_im;
  reg        [23:0]   shift_reg_32_re;
  reg        [23:0]   shift_reg_32_im;
  reg        [23:0]   shift_reg_33_re;
  reg        [23:0]   shift_reg_33_im;
  reg        [23:0]   shift_reg_34_re;
  reg        [23:0]   shift_reg_34_im;
  reg        [23:0]   shift_reg_35_re;
  reg        [23:0]   shift_reg_35_im;
  reg        [23:0]   shift_reg_36_re;
  reg        [23:0]   shift_reg_36_im;
  reg        [23:0]   shift_reg_37_re;
  reg        [23:0]   shift_reg_37_im;
  reg        [23:0]   shift_reg_38_re;
  reg        [23:0]   shift_reg_38_im;
  reg        [23:0]   shift_reg_39_re;
  reg        [23:0]   shift_reg_39_im;
  reg        [23:0]   shift_reg_40_re;
  reg        [23:0]   shift_reg_40_im;
  reg        [23:0]   shift_reg_41_re;
  reg        [23:0]   shift_reg_41_im;
  reg        [23:0]   shift_reg_42_re;
  reg        [23:0]   shift_reg_42_im;
  reg        [23:0]   shift_reg_43_re;
  reg        [23:0]   shift_reg_43_im;
  reg        [23:0]   shift_reg_44_re;
  reg        [23:0]   shift_reg_44_im;
  reg        [23:0]   shift_reg_45_re;
  reg        [23:0]   shift_reg_45_im;
  reg        [23:0]   shift_reg_46_re;
  reg        [23:0]   shift_reg_46_im;
  reg        [23:0]   shift_reg_47_re;
  reg        [23:0]   shift_reg_47_im;
  reg        [23:0]   shift_reg_48_re;
  reg        [23:0]   shift_reg_48_im;
  reg        [23:0]   shift_reg_49_re;
  reg        [23:0]   shift_reg_49_im;
  reg        [23:0]   shift_reg_50_re;
  reg        [23:0]   shift_reg_50_im;
  reg        [23:0]   shift_reg_51_re;
  reg        [23:0]   shift_reg_51_im;
  reg        [23:0]   shift_reg_52_re;
  reg        [23:0]   shift_reg_52_im;
  reg        [23:0]   shift_reg_53_re;
  reg        [23:0]   shift_reg_53_im;
  reg        [23:0]   shift_reg_54_re;
  reg        [23:0]   shift_reg_54_im;
  reg        [23:0]   shift_reg_55_re;
  reg        [23:0]   shift_reg_55_im;
  reg        [23:0]   shift_reg_56_re;
  reg        [23:0]   shift_reg_56_im;
  reg        [23:0]   shift_reg_57_re;
  reg        [23:0]   shift_reg_57_im;
  reg        [23:0]   shift_reg_58_re;
  reg        [23:0]   shift_reg_58_im;
  reg        [23:0]   shift_reg_59_re;
  reg        [23:0]   shift_reg_59_im;
  reg        [23:0]   shift_reg_60_re;
  reg        [23:0]   shift_reg_60_im;
  reg        [23:0]   shift_reg_61_re;
  reg        [23:0]   shift_reg_61_im;
  reg        [23:0]   shift_reg_62_re;
  reg        [23:0]   shift_reg_62_im;
  reg        [23:0]   shift_reg_63_re;
  reg        [23:0]   shift_reg_63_im;
  reg        [23:0]   shift_reg_64_re;
  reg        [23:0]   shift_reg_64_im;
  reg        [23:0]   shift_reg_65_re;
  reg        [23:0]   shift_reg_65_im;
  reg        [23:0]   shift_reg_66_re;
  reg        [23:0]   shift_reg_66_im;
  reg        [23:0]   shift_reg_67_re;
  reg        [23:0]   shift_reg_67_im;
  reg        [23:0]   shift_reg_68_re;
  reg        [23:0]   shift_reg_68_im;
  reg        [23:0]   shift_reg_69_re;
  reg        [23:0]   shift_reg_69_im;
  reg        [23:0]   shift_reg_70_re;
  reg        [23:0]   shift_reg_70_im;
  reg        [23:0]   shift_reg_71_re;
  reg        [23:0]   shift_reg_71_im;
  reg        [23:0]   shift_reg_72_re;
  reg        [23:0]   shift_reg_72_im;
  reg        [23:0]   shift_reg_73_re;
  reg        [23:0]   shift_reg_73_im;
  reg        [23:0]   shift_reg_74_re;
  reg        [23:0]   shift_reg_74_im;
  reg        [23:0]   shift_reg_75_re;
  reg        [23:0]   shift_reg_75_im;
  reg        [23:0]   shift_reg_76_re;
  reg        [23:0]   shift_reg_76_im;
  reg        [23:0]   shift_reg_77_re;
  reg        [23:0]   shift_reg_77_im;
  reg        [23:0]   shift_reg_78_re;
  reg        [23:0]   shift_reg_78_im;
  reg        [23:0]   shift_reg_79_re;
  reg        [23:0]   shift_reg_79_im;
  reg        [23:0]   shift_reg_80_re;
  reg        [23:0]   shift_reg_80_im;
  reg        [23:0]   shift_reg_81_re;
  reg        [23:0]   shift_reg_81_im;
  reg        [23:0]   shift_reg_82_re;
  reg        [23:0]   shift_reg_82_im;
  reg        [23:0]   shift_reg_83_re;
  reg        [23:0]   shift_reg_83_im;
  reg        [23:0]   shift_reg_84_re;
  reg        [23:0]   shift_reg_84_im;
  reg        [23:0]   shift_reg_85_re;
  reg        [23:0]   shift_reg_85_im;
  reg        [23:0]   shift_reg_86_re;
  reg        [23:0]   shift_reg_86_im;
  reg        [23:0]   shift_reg_87_re;
  reg        [23:0]   shift_reg_87_im;
  reg        [23:0]   shift_reg_88_re;
  reg        [23:0]   shift_reg_88_im;
  reg        [23:0]   shift_reg_89_re;
  reg        [23:0]   shift_reg_89_im;
  reg        [23:0]   shift_reg_90_re;
  reg        [23:0]   shift_reg_90_im;
  reg        [23:0]   shift_reg_91_re;
  reg        [23:0]   shift_reg_91_im;
  reg        [23:0]   shift_reg_92_re;
  reg        [23:0]   shift_reg_92_im;
  reg        [23:0]   shift_reg_93_re;
  reg        [23:0]   shift_reg_93_im;
  reg        [23:0]   shift_reg_94_re;
  reg        [23:0]   shift_reg_94_im;
  reg        [23:0]   shift_reg_95_re;
  reg        [23:0]   shift_reg_95_im;
  reg        [23:0]   shift_reg_96_re;
  reg        [23:0]   shift_reg_96_im;
  reg        [23:0]   shift_reg_97_re;
  reg        [23:0]   shift_reg_97_im;
  reg        [23:0]   shift_reg_98_re;
  reg        [23:0]   shift_reg_98_im;
  reg        [23:0]   shift_reg_99_re;
  reg        [23:0]   shift_reg_99_im;
  reg        [23:0]   shift_reg_100_re;
  reg        [23:0]   shift_reg_100_im;
  reg        [23:0]   shift_reg_101_re;
  reg        [23:0]   shift_reg_101_im;
  reg        [23:0]   shift_reg_102_re;
  reg        [23:0]   shift_reg_102_im;
  reg        [23:0]   shift_reg_103_re;
  reg        [23:0]   shift_reg_103_im;
  reg        [23:0]   shift_reg_104_re;
  reg        [23:0]   shift_reg_104_im;
  reg        [23:0]   shift_reg_105_re;
  reg        [23:0]   shift_reg_105_im;
  reg        [23:0]   shift_reg_106_re;
  reg        [23:0]   shift_reg_106_im;
  reg        [23:0]   shift_reg_107_re;
  reg        [23:0]   shift_reg_107_im;
  reg        [23:0]   shift_reg_108_re;
  reg        [23:0]   shift_reg_108_im;
  reg        [23:0]   shift_reg_109_re;
  reg        [23:0]   shift_reg_109_im;
  reg        [23:0]   shift_reg_110_re;
  reg        [23:0]   shift_reg_110_im;
  reg        [23:0]   shift_reg_111_re;
  reg        [23:0]   shift_reg_111_im;
  reg        [23:0]   shift_reg_112_re;
  reg        [23:0]   shift_reg_112_im;
  reg        [23:0]   shift_reg_113_re;
  reg        [23:0]   shift_reg_113_im;
  reg        [23:0]   shift_reg_114_re;
  reg        [23:0]   shift_reg_114_im;
  reg        [23:0]   shift_reg_115_re;
  reg        [23:0]   shift_reg_115_im;
  reg        [23:0]   shift_reg_116_re;
  reg        [23:0]   shift_reg_116_im;
  reg        [23:0]   shift_reg_117_re;
  reg        [23:0]   shift_reg_117_im;
  reg        [23:0]   shift_reg_118_re;
  reg        [23:0]   shift_reg_118_im;
  reg        [23:0]   shift_reg_119_re;
  reg        [23:0]   shift_reg_119_im;
  reg        [23:0]   shift_reg_120_re;
  reg        [23:0]   shift_reg_120_im;
  reg        [23:0]   shift_reg_121_re;
  reg        [23:0]   shift_reg_121_im;
  reg        [23:0]   shift_reg_122_re;
  reg        [23:0]   shift_reg_122_im;
  reg        [23:0]   shift_reg_123_re;
  reg        [23:0]   shift_reg_123_im;
  reg        [23:0]   shift_reg_124_re;
  reg        [23:0]   shift_reg_124_im;
  reg        [23:0]   shift_reg_125_re;
  reg        [23:0]   shift_reg_125_im;
  reg        [23:0]   shift_reg_126_re;
  reg        [23:0]   shift_reg_126_im;
  reg        [23:0]   shift_reg_127_re;
  reg        [23:0]   shift_reg_127_im;
  reg        [23:0]   shift_reg_128_re;
  reg        [23:0]   shift_reg_128_im;
  reg        [23:0]   shift_reg_129_re;
  reg        [23:0]   shift_reg_129_im;
  reg        [23:0]   shift_reg_130_re;
  reg        [23:0]   shift_reg_130_im;
  reg        [23:0]   shift_reg_131_re;
  reg        [23:0]   shift_reg_131_im;
  reg        [23:0]   shift_reg_132_re;
  reg        [23:0]   shift_reg_132_im;
  reg        [23:0]   shift_reg_133_re;
  reg        [23:0]   shift_reg_133_im;
  reg        [23:0]   shift_reg_134_re;
  reg        [23:0]   shift_reg_134_im;
  reg        [23:0]   shift_reg_135_re;
  reg        [23:0]   shift_reg_135_im;
  reg        [23:0]   shift_reg_136_re;
  reg        [23:0]   shift_reg_136_im;
  reg        [23:0]   shift_reg_137_re;
  reg        [23:0]   shift_reg_137_im;
  reg        [23:0]   shift_reg_138_re;
  reg        [23:0]   shift_reg_138_im;
  reg        [23:0]   shift_reg_139_re;
  reg        [23:0]   shift_reg_139_im;
  reg        [23:0]   shift_reg_140_re;
  reg        [23:0]   shift_reg_140_im;
  reg        [23:0]   shift_reg_141_re;
  reg        [23:0]   shift_reg_141_im;
  reg        [23:0]   shift_reg_142_re;
  reg        [23:0]   shift_reg_142_im;
  reg        [23:0]   shift_reg_143_re;
  reg        [23:0]   shift_reg_143_im;
  reg        [23:0]   shift_reg_144_re;
  reg        [23:0]   shift_reg_144_im;
  reg        [23:0]   shift_reg_145_re;
  reg        [23:0]   shift_reg_145_im;
  reg        [23:0]   shift_reg_146_re;
  reg        [23:0]   shift_reg_146_im;
  reg        [23:0]   shift_reg_147_re;
  reg        [23:0]   shift_reg_147_im;
  reg        [23:0]   shift_reg_148_re;
  reg        [23:0]   shift_reg_148_im;
  reg        [23:0]   shift_reg_149_re;
  reg        [23:0]   shift_reg_149_im;
  reg        [23:0]   shift_reg_150_re;
  reg        [23:0]   shift_reg_150_im;
  reg        [23:0]   shift_reg_151_re;
  reg        [23:0]   shift_reg_151_im;
  reg        [23:0]   shift_reg_152_re;
  reg        [23:0]   shift_reg_152_im;
  reg        [23:0]   shift_reg_153_re;
  reg        [23:0]   shift_reg_153_im;
  reg        [23:0]   shift_reg_154_re;
  reg        [23:0]   shift_reg_154_im;
  reg        [23:0]   shift_reg_155_re;
  reg        [23:0]   shift_reg_155_im;
  reg        [23:0]   shift_reg_156_re;
  reg        [23:0]   shift_reg_156_im;
  reg        [23:0]   shift_reg_157_re;
  reg        [23:0]   shift_reg_157_im;
  reg        [23:0]   shift_reg_158_re;
  reg        [23:0]   shift_reg_158_im;
  reg        [23:0]   shift_reg_159_re;
  reg        [23:0]   shift_reg_159_im;
  reg        [23:0]   shift_reg_160_re;
  reg        [23:0]   shift_reg_160_im;
  reg        [23:0]   shift_reg_161_re;
  reg        [23:0]   shift_reg_161_im;
  reg        [23:0]   shift_reg_162_re;
  reg        [23:0]   shift_reg_162_im;
  reg        [23:0]   shift_reg_163_re;
  reg        [23:0]   shift_reg_163_im;
  reg        [23:0]   shift_reg_164_re;
  reg        [23:0]   shift_reg_164_im;
  reg        [23:0]   shift_reg_165_re;
  reg        [23:0]   shift_reg_165_im;
  reg        [23:0]   shift_reg_166_re;
  reg        [23:0]   shift_reg_166_im;
  reg        [23:0]   shift_reg_167_re;
  reg        [23:0]   shift_reg_167_im;
  reg        [23:0]   shift_reg_168_re;
  reg        [23:0]   shift_reg_168_im;
  reg        [23:0]   shift_reg_169_re;
  reg        [23:0]   shift_reg_169_im;
  reg        [23:0]   shift_reg_170_re;
  reg        [23:0]   shift_reg_170_im;
  reg        [23:0]   shift_reg_171_re;
  reg        [23:0]   shift_reg_171_im;
  reg        [23:0]   shift_reg_172_re;
  reg        [23:0]   shift_reg_172_im;
  reg        [23:0]   shift_reg_173_re;
  reg        [23:0]   shift_reg_173_im;
  reg        [23:0]   shift_reg_174_re;
  reg        [23:0]   shift_reg_174_im;
  reg        [23:0]   shift_reg_175_re;
  reg        [23:0]   shift_reg_175_im;
  reg        [23:0]   shift_reg_176_re;
  reg        [23:0]   shift_reg_176_im;
  reg        [23:0]   shift_reg_177_re;
  reg        [23:0]   shift_reg_177_im;
  reg        [23:0]   shift_reg_178_re;
  reg        [23:0]   shift_reg_178_im;
  reg        [23:0]   shift_reg_179_re;
  reg        [23:0]   shift_reg_179_im;
  reg        [23:0]   shift_reg_180_re;
  reg        [23:0]   shift_reg_180_im;
  reg        [23:0]   shift_reg_181_re;
  reg        [23:0]   shift_reg_181_im;
  reg        [23:0]   shift_reg_182_re;
  reg        [23:0]   shift_reg_182_im;
  reg        [23:0]   shift_reg_183_re;
  reg        [23:0]   shift_reg_183_im;
  reg        [23:0]   shift_reg_184_re;
  reg        [23:0]   shift_reg_184_im;
  reg        [23:0]   shift_reg_185_re;
  reg        [23:0]   shift_reg_185_im;
  reg        [23:0]   shift_reg_186_re;
  reg        [23:0]   shift_reg_186_im;
  reg        [23:0]   shift_reg_187_re;
  reg        [23:0]   shift_reg_187_im;
  reg        [23:0]   shift_reg_188_re;
  reg        [23:0]   shift_reg_188_im;
  reg        [23:0]   shift_reg_189_re;
  reg        [23:0]   shift_reg_189_im;
  reg        [23:0]   shift_reg_190_re;
  reg        [23:0]   shift_reg_190_im;
  reg        [23:0]   shift_reg_191_re;
  reg        [23:0]   shift_reg_191_im;
  reg        [23:0]   shift_reg_192_re;
  reg        [23:0]   shift_reg_192_im;
  reg        [23:0]   shift_reg_193_re;
  reg        [23:0]   shift_reg_193_im;
  reg        [23:0]   shift_reg_194_re;
  reg        [23:0]   shift_reg_194_im;
  reg        [23:0]   shift_reg_195_re;
  reg        [23:0]   shift_reg_195_im;
  reg        [23:0]   shift_reg_196_re;
  reg        [23:0]   shift_reg_196_im;
  reg        [23:0]   shift_reg_197_re;
  reg        [23:0]   shift_reg_197_im;
  reg        [23:0]   shift_reg_198_re;
  reg        [23:0]   shift_reg_198_im;
  reg        [23:0]   shift_reg_199_re;
  reg        [23:0]   shift_reg_199_im;
  reg        [23:0]   shift_reg_200_re;
  reg        [23:0]   shift_reg_200_im;
  reg        [23:0]   shift_reg_201_re;
  reg        [23:0]   shift_reg_201_im;
  reg        [23:0]   shift_reg_202_re;
  reg        [23:0]   shift_reg_202_im;
  reg        [23:0]   shift_reg_203_re;
  reg        [23:0]   shift_reg_203_im;
  reg        [23:0]   shift_reg_204_re;
  reg        [23:0]   shift_reg_204_im;
  reg        [23:0]   shift_reg_205_re;
  reg        [23:0]   shift_reg_205_im;
  reg        [23:0]   shift_reg_206_re;
  reg        [23:0]   shift_reg_206_im;
  reg        [23:0]   shift_reg_207_re;
  reg        [23:0]   shift_reg_207_im;
  reg        [23:0]   shift_reg_208_re;
  reg        [23:0]   shift_reg_208_im;
  reg        [23:0]   shift_reg_209_re;
  reg        [23:0]   shift_reg_209_im;
  reg        [23:0]   shift_reg_210_re;
  reg        [23:0]   shift_reg_210_im;
  reg        [23:0]   shift_reg_211_re;
  reg        [23:0]   shift_reg_211_im;
  reg        [23:0]   shift_reg_212_re;
  reg        [23:0]   shift_reg_212_im;
  reg        [23:0]   shift_reg_213_re;
  reg        [23:0]   shift_reg_213_im;
  reg        [23:0]   shift_reg_214_re;
  reg        [23:0]   shift_reg_214_im;
  reg        [23:0]   shift_reg_215_re;
  reg        [23:0]   shift_reg_215_im;
  reg        [23:0]   shift_reg_216_re;
  reg        [23:0]   shift_reg_216_im;
  reg        [23:0]   shift_reg_217_re;
  reg        [23:0]   shift_reg_217_im;
  reg        [23:0]   shift_reg_218_re;
  reg        [23:0]   shift_reg_218_im;
  reg        [23:0]   shift_reg_219_re;
  reg        [23:0]   shift_reg_219_im;
  reg        [23:0]   shift_reg_220_re;
  reg        [23:0]   shift_reg_220_im;
  reg        [23:0]   shift_reg_221_re;
  reg        [23:0]   shift_reg_221_im;
  reg        [23:0]   shift_reg_222_re;
  reg        [23:0]   shift_reg_222_im;
  reg        [23:0]   shift_reg_223_re;
  reg        [23:0]   shift_reg_223_im;
  reg        [23:0]   shift_reg_224_re;
  reg        [23:0]   shift_reg_224_im;
  reg        [23:0]   shift_reg_225_re;
  reg        [23:0]   shift_reg_225_im;
  reg        [23:0]   shift_reg_226_re;
  reg        [23:0]   shift_reg_226_im;
  reg        [23:0]   shift_reg_227_re;
  reg        [23:0]   shift_reg_227_im;
  reg        [23:0]   shift_reg_228_re;
  reg        [23:0]   shift_reg_228_im;
  reg        [23:0]   shift_reg_229_re;
  reg        [23:0]   shift_reg_229_im;
  reg        [23:0]   shift_reg_230_re;
  reg        [23:0]   shift_reg_230_im;
  reg        [23:0]   shift_reg_231_re;
  reg        [23:0]   shift_reg_231_im;
  reg        [23:0]   shift_reg_232_re;
  reg        [23:0]   shift_reg_232_im;
  reg        [23:0]   shift_reg_233_re;
  reg        [23:0]   shift_reg_233_im;
  reg        [23:0]   shift_reg_234_re;
  reg        [23:0]   shift_reg_234_im;
  reg        [23:0]   shift_reg_235_re;
  reg        [23:0]   shift_reg_235_im;
  reg        [23:0]   shift_reg_236_re;
  reg        [23:0]   shift_reg_236_im;
  reg        [23:0]   shift_reg_237_re;
  reg        [23:0]   shift_reg_237_im;
  reg        [23:0]   shift_reg_238_re;
  reg        [23:0]   shift_reg_238_im;
  reg        [23:0]   shift_reg_239_re;
  reg        [23:0]   shift_reg_239_im;
  reg        [23:0]   shift_reg_240_re;
  reg        [23:0]   shift_reg_240_im;
  reg        [23:0]   shift_reg_241_re;
  reg        [23:0]   shift_reg_241_im;
  reg        [23:0]   shift_reg_242_re;
  reg        [23:0]   shift_reg_242_im;
  reg        [23:0]   shift_reg_243_re;
  reg        [23:0]   shift_reg_243_im;
  reg        [23:0]   shift_reg_244_re;
  reg        [23:0]   shift_reg_244_im;
  reg        [23:0]   shift_reg_245_re;
  reg        [23:0]   shift_reg_245_im;
  reg        [23:0]   shift_reg_246_re;
  reg        [23:0]   shift_reg_246_im;
  reg        [23:0]   shift_reg_247_re;
  reg        [23:0]   shift_reg_247_im;
  reg        [23:0]   shift_reg_248_re;
  reg        [23:0]   shift_reg_248_im;
  reg        [23:0]   shift_reg_249_re;
  reg        [23:0]   shift_reg_249_im;
  reg        [23:0]   shift_reg_250_re;
  reg        [23:0]   shift_reg_250_im;
  reg        [23:0]   shift_reg_251_re;
  reg        [23:0]   shift_reg_251_im;
  reg        [23:0]   shift_reg_252_re;
  reg        [23:0]   shift_reg_252_im;
  reg        [23:0]   shift_reg_253_re;
  reg        [23:0]   shift_reg_253_im;
  reg        [23:0]   shift_reg_254_re;
  reg        [23:0]   shift_reg_254_im;
  reg        [23:0]   shift_reg_255_re;
  reg        [23:0]   shift_reg_255_im;
  reg        [23:0]   shift_reg_256_re;
  reg        [23:0]   shift_reg_256_im;
  reg        [23:0]   shift_reg_257_re;
  reg        [23:0]   shift_reg_257_im;
  reg        [23:0]   shift_reg_258_re;
  reg        [23:0]   shift_reg_258_im;
  reg        [23:0]   shift_reg_259_re;
  reg        [23:0]   shift_reg_259_im;
  reg        [23:0]   shift_reg_260_re;
  reg        [23:0]   shift_reg_260_im;
  reg        [23:0]   shift_reg_261_re;
  reg        [23:0]   shift_reg_261_im;
  reg        [23:0]   shift_reg_262_re;
  reg        [23:0]   shift_reg_262_im;
  reg        [23:0]   shift_reg_263_re;
  reg        [23:0]   shift_reg_263_im;
  reg        [23:0]   shift_reg_264_re;
  reg        [23:0]   shift_reg_264_im;
  reg        [23:0]   shift_reg_265_re;
  reg        [23:0]   shift_reg_265_im;
  reg        [23:0]   shift_reg_266_re;
  reg        [23:0]   shift_reg_266_im;
  reg        [23:0]   shift_reg_267_re;
  reg        [23:0]   shift_reg_267_im;
  reg        [23:0]   shift_reg_268_re;
  reg        [23:0]   shift_reg_268_im;
  reg        [23:0]   shift_reg_269_re;
  reg        [23:0]   shift_reg_269_im;
  reg        [23:0]   shift_reg_270_re;
  reg        [23:0]   shift_reg_270_im;
  reg        [23:0]   shift_reg_271_re;
  reg        [23:0]   shift_reg_271_im;
  reg        [23:0]   shift_reg_272_re;
  reg        [23:0]   shift_reg_272_im;
  reg        [23:0]   shift_reg_273_re;
  reg        [23:0]   shift_reg_273_im;
  reg        [23:0]   shift_reg_274_re;
  reg        [23:0]   shift_reg_274_im;
  reg        [23:0]   shift_reg_275_re;
  reg        [23:0]   shift_reg_275_im;
  reg        [23:0]   shift_reg_276_re;
  reg        [23:0]   shift_reg_276_im;
  reg        [23:0]   shift_reg_277_re;
  reg        [23:0]   shift_reg_277_im;
  reg        [23:0]   shift_reg_278_re;
  reg        [23:0]   shift_reg_278_im;
  reg        [23:0]   shift_reg_279_re;
  reg        [23:0]   shift_reg_279_im;
  reg        [23:0]   shift_reg_280_re;
  reg        [23:0]   shift_reg_280_im;
  reg        [23:0]   shift_reg_281_re;
  reg        [23:0]   shift_reg_281_im;
  reg        [23:0]   shift_reg_282_re;
  reg        [23:0]   shift_reg_282_im;
  reg        [23:0]   shift_reg_283_re;
  reg        [23:0]   shift_reg_283_im;
  reg        [23:0]   shift_reg_284_re;
  reg        [23:0]   shift_reg_284_im;
  reg        [23:0]   shift_reg_285_re;
  reg        [23:0]   shift_reg_285_im;
  reg        [23:0]   shift_reg_286_re;
  reg        [23:0]   shift_reg_286_im;
  reg        [23:0]   shift_reg_287_re;
  reg        [23:0]   shift_reg_287_im;
  reg        [23:0]   shift_reg_288_re;
  reg        [23:0]   shift_reg_288_im;
  reg        [23:0]   shift_reg_289_re;
  reg        [23:0]   shift_reg_289_im;
  reg        [23:0]   shift_reg_290_re;
  reg        [23:0]   shift_reg_290_im;
  reg        [23:0]   shift_reg_291_re;
  reg        [23:0]   shift_reg_291_im;
  reg        [23:0]   shift_reg_292_re;
  reg        [23:0]   shift_reg_292_im;
  reg        [23:0]   shift_reg_293_re;
  reg        [23:0]   shift_reg_293_im;
  reg        [23:0]   shift_reg_294_re;
  reg        [23:0]   shift_reg_294_im;
  reg        [23:0]   shift_reg_295_re;
  reg        [23:0]   shift_reg_295_im;
  reg        [23:0]   shift_reg_296_re;
  reg        [23:0]   shift_reg_296_im;
  reg        [23:0]   shift_reg_297_re;
  reg        [23:0]   shift_reg_297_im;
  reg        [23:0]   shift_reg_298_re;
  reg        [23:0]   shift_reg_298_im;
  reg        [23:0]   shift_reg_299_re;
  reg        [23:0]   shift_reg_299_im;
  reg        [23:0]   shift_reg_300_re;
  reg        [23:0]   shift_reg_300_im;
  reg        [23:0]   shift_reg_301_re;
  reg        [23:0]   shift_reg_301_im;
  reg        [23:0]   shift_reg_302_re;
  reg        [23:0]   shift_reg_302_im;
  reg        [23:0]   shift_reg_303_re;
  reg        [23:0]   shift_reg_303_im;
  reg        [23:0]   shift_reg_304_re;
  reg        [23:0]   shift_reg_304_im;
  reg        [23:0]   shift_reg_305_re;
  reg        [23:0]   shift_reg_305_im;
  reg        [23:0]   shift_reg_306_re;
  reg        [23:0]   shift_reg_306_im;
  reg        [23:0]   shift_reg_307_re;
  reg        [23:0]   shift_reg_307_im;
  reg        [23:0]   shift_reg_308_re;
  reg        [23:0]   shift_reg_308_im;
  reg        [23:0]   shift_reg_309_re;
  reg        [23:0]   shift_reg_309_im;
  reg        [23:0]   shift_reg_310_re;
  reg        [23:0]   shift_reg_310_im;
  reg        [23:0]   shift_reg_311_re;
  reg        [23:0]   shift_reg_311_im;
  reg        [23:0]   shift_reg_312_re;
  reg        [23:0]   shift_reg_312_im;
  reg        [23:0]   shift_reg_313_re;
  reg        [23:0]   shift_reg_313_im;
  reg        [23:0]   shift_reg_314_re;
  reg        [23:0]   shift_reg_314_im;
  reg        [23:0]   shift_reg_315_re;
  reg        [23:0]   shift_reg_315_im;
  reg        [23:0]   shift_reg_316_re;
  reg        [23:0]   shift_reg_316_im;
  reg        [23:0]   shift_reg_317_re;
  reg        [23:0]   shift_reg_317_im;
  reg        [23:0]   shift_reg_318_re;
  reg        [23:0]   shift_reg_318_im;
  reg        [23:0]   shift_reg_319_re;
  reg        [23:0]   shift_reg_319_im;
  reg        [23:0]   shift_reg_320_re;
  reg        [23:0]   shift_reg_320_im;
  reg        [23:0]   shift_reg_321_re;
  reg        [23:0]   shift_reg_321_im;
  reg        [23:0]   shift_reg_322_re;
  reg        [23:0]   shift_reg_322_im;
  reg        [23:0]   shift_reg_323_re;
  reg        [23:0]   shift_reg_323_im;
  reg        [23:0]   shift_reg_324_re;
  reg        [23:0]   shift_reg_324_im;
  reg        [23:0]   shift_reg_325_re;
  reg        [23:0]   shift_reg_325_im;
  reg        [23:0]   shift_reg_326_re;
  reg        [23:0]   shift_reg_326_im;
  reg        [23:0]   shift_reg_327_re;
  reg        [23:0]   shift_reg_327_im;
  reg        [23:0]   shift_reg_328_re;
  reg        [23:0]   shift_reg_328_im;
  reg        [23:0]   shift_reg_329_re;
  reg        [23:0]   shift_reg_329_im;
  reg        [23:0]   shift_reg_330_re;
  reg        [23:0]   shift_reg_330_im;
  reg        [23:0]   shift_reg_331_re;
  reg        [23:0]   shift_reg_331_im;
  reg        [23:0]   shift_reg_332_re;
  reg        [23:0]   shift_reg_332_im;
  reg        [23:0]   shift_reg_333_re;
  reg        [23:0]   shift_reg_333_im;
  reg        [23:0]   shift_reg_334_re;
  reg        [23:0]   shift_reg_334_im;
  reg        [23:0]   shift_reg_335_re;
  reg        [23:0]   shift_reg_335_im;
  reg        [23:0]   shift_reg_336_re;
  reg        [23:0]   shift_reg_336_im;
  reg        [23:0]   shift_reg_337_re;
  reg        [23:0]   shift_reg_337_im;
  reg        [23:0]   shift_reg_338_re;
  reg        [23:0]   shift_reg_338_im;
  reg        [23:0]   shift_reg_339_re;
  reg        [23:0]   shift_reg_339_im;
  reg        [23:0]   shift_reg_340_re;
  reg        [23:0]   shift_reg_340_im;
  reg        [23:0]   shift_reg_341_re;
  reg        [23:0]   shift_reg_341_im;
  reg        [23:0]   shift_reg_342_re;
  reg        [23:0]   shift_reg_342_im;
  reg        [23:0]   shift_reg_343_re;
  reg        [23:0]   shift_reg_343_im;
  reg        [23:0]   shift_reg_344_re;
  reg        [23:0]   shift_reg_344_im;
  reg        [23:0]   shift_reg_345_re;
  reg        [23:0]   shift_reg_345_im;
  reg        [23:0]   shift_reg_346_re;
  reg        [23:0]   shift_reg_346_im;
  reg        [23:0]   shift_reg_347_re;
  reg        [23:0]   shift_reg_347_im;
  reg        [23:0]   shift_reg_348_re;
  reg        [23:0]   shift_reg_348_im;
  reg        [23:0]   shift_reg_349_re;
  reg        [23:0]   shift_reg_349_im;
  reg        [23:0]   shift_reg_350_re;
  reg        [23:0]   shift_reg_350_im;
  reg        [23:0]   shift_reg_351_re;
  reg        [23:0]   shift_reg_351_im;
  reg        [23:0]   shift_reg_352_re;
  reg        [23:0]   shift_reg_352_im;
  reg        [23:0]   shift_reg_353_re;
  reg        [23:0]   shift_reg_353_im;
  reg        [23:0]   shift_reg_354_re;
  reg        [23:0]   shift_reg_354_im;
  reg        [23:0]   shift_reg_355_re;
  reg        [23:0]   shift_reg_355_im;
  reg        [23:0]   shift_reg_356_re;
  reg        [23:0]   shift_reg_356_im;
  reg        [23:0]   shift_reg_357_re;
  reg        [23:0]   shift_reg_357_im;
  reg        [23:0]   shift_reg_358_re;
  reg        [23:0]   shift_reg_358_im;
  reg        [23:0]   shift_reg_359_re;
  reg        [23:0]   shift_reg_359_im;
  reg        [23:0]   shift_reg_360_re;
  reg        [23:0]   shift_reg_360_im;
  reg        [23:0]   shift_reg_361_re;
  reg        [23:0]   shift_reg_361_im;
  reg        [23:0]   shift_reg_362_re;
  reg        [23:0]   shift_reg_362_im;
  reg        [23:0]   shift_reg_363_re;
  reg        [23:0]   shift_reg_363_im;
  reg        [23:0]   shift_reg_364_re;
  reg        [23:0]   shift_reg_364_im;
  reg        [23:0]   shift_reg_365_re;
  reg        [23:0]   shift_reg_365_im;
  reg        [23:0]   shift_reg_366_re;
  reg        [23:0]   shift_reg_366_im;
  reg        [23:0]   shift_reg_367_re;
  reg        [23:0]   shift_reg_367_im;
  reg        [23:0]   shift_reg_368_re;
  reg        [23:0]   shift_reg_368_im;
  reg        [23:0]   shift_reg_369_re;
  reg        [23:0]   shift_reg_369_im;
  reg        [23:0]   shift_reg_370_re;
  reg        [23:0]   shift_reg_370_im;
  reg        [23:0]   shift_reg_371_re;
  reg        [23:0]   shift_reg_371_im;
  reg        [23:0]   shift_reg_372_re;
  reg        [23:0]   shift_reg_372_im;
  reg        [23:0]   shift_reg_373_re;
  reg        [23:0]   shift_reg_373_im;
  reg        [23:0]   shift_reg_374_re;
  reg        [23:0]   shift_reg_374_im;
  reg        [23:0]   shift_reg_375_re;
  reg        [23:0]   shift_reg_375_im;
  reg        [23:0]   shift_reg_376_re;
  reg        [23:0]   shift_reg_376_im;
  reg        [23:0]   shift_reg_377_re;
  reg        [23:0]   shift_reg_377_im;
  reg        [23:0]   shift_reg_378_re;
  reg        [23:0]   shift_reg_378_im;
  reg        [23:0]   shift_reg_379_re;
  reg        [23:0]   shift_reg_379_im;
  reg        [23:0]   shift_reg_380_re;
  reg        [23:0]   shift_reg_380_im;
  reg        [23:0]   shift_reg_381_re;
  reg        [23:0]   shift_reg_381_im;
  reg        [23:0]   shift_reg_382_re;
  reg        [23:0]   shift_reg_382_im;
  reg        [23:0]   shift_reg_383_re;
  reg        [23:0]   shift_reg_383_im;
  reg        [23:0]   shift_reg_384_re;
  reg        [23:0]   shift_reg_384_im;
  reg        [23:0]   shift_reg_385_re;
  reg        [23:0]   shift_reg_385_im;
  reg        [23:0]   shift_reg_386_re;
  reg        [23:0]   shift_reg_386_im;
  reg        [23:0]   shift_reg_387_re;
  reg        [23:0]   shift_reg_387_im;
  reg        [23:0]   shift_reg_388_re;
  reg        [23:0]   shift_reg_388_im;
  reg        [23:0]   shift_reg_389_re;
  reg        [23:0]   shift_reg_389_im;
  reg        [23:0]   shift_reg_390_re;
  reg        [23:0]   shift_reg_390_im;
  reg        [23:0]   shift_reg_391_re;
  reg        [23:0]   shift_reg_391_im;
  reg        [23:0]   shift_reg_392_re;
  reg        [23:0]   shift_reg_392_im;
  reg        [23:0]   shift_reg_393_re;
  reg        [23:0]   shift_reg_393_im;
  reg        [23:0]   shift_reg_394_re;
  reg        [23:0]   shift_reg_394_im;
  reg        [23:0]   shift_reg_395_re;
  reg        [23:0]   shift_reg_395_im;
  reg        [23:0]   shift_reg_396_re;
  reg        [23:0]   shift_reg_396_im;
  reg        [23:0]   shift_reg_397_re;
  reg        [23:0]   shift_reg_397_im;
  reg        [23:0]   shift_reg_398_re;
  reg        [23:0]   shift_reg_398_im;
  reg        [23:0]   shift_reg_399_re;
  reg        [23:0]   shift_reg_399_im;
  reg        [23:0]   shift_reg_400_re;
  reg        [23:0]   shift_reg_400_im;
  reg        [23:0]   shift_reg_401_re;
  reg        [23:0]   shift_reg_401_im;
  reg        [23:0]   shift_reg_402_re;
  reg        [23:0]   shift_reg_402_im;
  reg        [23:0]   shift_reg_403_re;
  reg        [23:0]   shift_reg_403_im;
  reg        [23:0]   shift_reg_404_re;
  reg        [23:0]   shift_reg_404_im;
  reg        [23:0]   shift_reg_405_re;
  reg        [23:0]   shift_reg_405_im;
  reg        [23:0]   shift_reg_406_re;
  reg        [23:0]   shift_reg_406_im;
  reg        [23:0]   shift_reg_407_re;
  reg        [23:0]   shift_reg_407_im;
  reg        [23:0]   shift_reg_408_re;
  reg        [23:0]   shift_reg_408_im;
  reg        [23:0]   shift_reg_409_re;
  reg        [23:0]   shift_reg_409_im;
  reg        [23:0]   shift_reg_410_re;
  reg        [23:0]   shift_reg_410_im;
  reg        [23:0]   shift_reg_411_re;
  reg        [23:0]   shift_reg_411_im;
  reg        [23:0]   shift_reg_412_re;
  reg        [23:0]   shift_reg_412_im;
  reg        [23:0]   shift_reg_413_re;
  reg        [23:0]   shift_reg_413_im;
  reg        [23:0]   shift_reg_414_re;
  reg        [23:0]   shift_reg_414_im;
  reg        [23:0]   shift_reg_415_re;
  reg        [23:0]   shift_reg_415_im;
  reg        [23:0]   shift_reg_416_re;
  reg        [23:0]   shift_reg_416_im;
  reg        [23:0]   shift_reg_417_re;
  reg        [23:0]   shift_reg_417_im;
  reg        [23:0]   shift_reg_418_re;
  reg        [23:0]   shift_reg_418_im;
  reg        [23:0]   shift_reg_419_re;
  reg        [23:0]   shift_reg_419_im;
  reg        [23:0]   shift_reg_420_re;
  reg        [23:0]   shift_reg_420_im;
  reg        [23:0]   shift_reg_421_re;
  reg        [23:0]   shift_reg_421_im;
  reg        [23:0]   shift_reg_422_re;
  reg        [23:0]   shift_reg_422_im;
  reg        [23:0]   shift_reg_423_re;
  reg        [23:0]   shift_reg_423_im;
  reg        [23:0]   shift_reg_424_re;
  reg        [23:0]   shift_reg_424_im;
  reg        [23:0]   shift_reg_425_re;
  reg        [23:0]   shift_reg_425_im;
  reg        [23:0]   shift_reg_426_re;
  reg        [23:0]   shift_reg_426_im;
  reg        [23:0]   shift_reg_427_re;
  reg        [23:0]   shift_reg_427_im;
  reg        [23:0]   shift_reg_428_re;
  reg        [23:0]   shift_reg_428_im;
  reg        [23:0]   shift_reg_429_re;
  reg        [23:0]   shift_reg_429_im;
  reg        [23:0]   shift_reg_430_re;
  reg        [23:0]   shift_reg_430_im;
  reg        [23:0]   shift_reg_431_re;
  reg        [23:0]   shift_reg_431_im;
  reg        [23:0]   shift_reg_432_re;
  reg        [23:0]   shift_reg_432_im;
  reg        [23:0]   shift_reg_433_re;
  reg        [23:0]   shift_reg_433_im;
  reg        [23:0]   shift_reg_434_re;
  reg        [23:0]   shift_reg_434_im;
  reg        [23:0]   shift_reg_435_re;
  reg        [23:0]   shift_reg_435_im;
  reg        [23:0]   shift_reg_436_re;
  reg        [23:0]   shift_reg_436_im;
  reg        [23:0]   shift_reg_437_re;
  reg        [23:0]   shift_reg_437_im;
  reg        [23:0]   shift_reg_438_re;
  reg        [23:0]   shift_reg_438_im;
  reg        [23:0]   shift_reg_439_re;
  reg        [23:0]   shift_reg_439_im;
  reg        [23:0]   shift_reg_440_re;
  reg        [23:0]   shift_reg_440_im;
  reg        [23:0]   shift_reg_441_re;
  reg        [23:0]   shift_reg_441_im;
  reg        [23:0]   shift_reg_442_re;
  reg        [23:0]   shift_reg_442_im;
  reg        [23:0]   shift_reg_443_re;
  reg        [23:0]   shift_reg_443_im;
  reg        [23:0]   shift_reg_444_re;
  reg        [23:0]   shift_reg_444_im;
  reg        [23:0]   shift_reg_445_re;
  reg        [23:0]   shift_reg_445_im;
  reg        [23:0]   shift_reg_446_re;
  reg        [23:0]   shift_reg_446_im;
  reg        [23:0]   shift_reg_447_re;
  reg        [23:0]   shift_reg_447_im;
  reg        [23:0]   shift_reg_448_re;
  reg        [23:0]   shift_reg_448_im;
  reg        [23:0]   shift_reg_449_re;
  reg        [23:0]   shift_reg_449_im;
  reg        [23:0]   shift_reg_450_re;
  reg        [23:0]   shift_reg_450_im;
  reg        [23:0]   shift_reg_451_re;
  reg        [23:0]   shift_reg_451_im;
  reg        [23:0]   shift_reg_452_re;
  reg        [23:0]   shift_reg_452_im;
  reg        [23:0]   shift_reg_453_re;
  reg        [23:0]   shift_reg_453_im;
  reg        [23:0]   shift_reg_454_re;
  reg        [23:0]   shift_reg_454_im;
  reg        [23:0]   shift_reg_455_re;
  reg        [23:0]   shift_reg_455_im;
  reg        [23:0]   shift_reg_456_re;
  reg        [23:0]   shift_reg_456_im;
  reg        [23:0]   shift_reg_457_re;
  reg        [23:0]   shift_reg_457_im;
  reg        [23:0]   shift_reg_458_re;
  reg        [23:0]   shift_reg_458_im;
  reg        [23:0]   shift_reg_459_re;
  reg        [23:0]   shift_reg_459_im;
  reg        [23:0]   shift_reg_460_re;
  reg        [23:0]   shift_reg_460_im;
  reg        [23:0]   shift_reg_461_re;
  reg        [23:0]   shift_reg_461_im;
  reg        [23:0]   shift_reg_462_re;
  reg        [23:0]   shift_reg_462_im;
  reg        [23:0]   shift_reg_463_re;
  reg        [23:0]   shift_reg_463_im;
  reg        [23:0]   shift_reg_464_re;
  reg        [23:0]   shift_reg_464_im;
  reg        [23:0]   shift_reg_465_re;
  reg        [23:0]   shift_reg_465_im;
  reg        [23:0]   shift_reg_466_re;
  reg        [23:0]   shift_reg_466_im;
  reg        [23:0]   shift_reg_467_re;
  reg        [23:0]   shift_reg_467_im;
  reg        [23:0]   shift_reg_468_re;
  reg        [23:0]   shift_reg_468_im;
  reg        [23:0]   shift_reg_469_re;
  reg        [23:0]   shift_reg_469_im;
  reg        [23:0]   shift_reg_470_re;
  reg        [23:0]   shift_reg_470_im;
  reg        [23:0]   shift_reg_471_re;
  reg        [23:0]   shift_reg_471_im;
  reg        [23:0]   shift_reg_472_re;
  reg        [23:0]   shift_reg_472_im;
  reg        [23:0]   shift_reg_473_re;
  reg        [23:0]   shift_reg_473_im;
  reg        [23:0]   shift_reg_474_re;
  reg        [23:0]   shift_reg_474_im;
  reg        [23:0]   shift_reg_475_re;
  reg        [23:0]   shift_reg_475_im;
  reg        [23:0]   shift_reg_476_re;
  reg        [23:0]   shift_reg_476_im;
  reg        [23:0]   shift_reg_477_re;
  reg        [23:0]   shift_reg_477_im;
  reg        [23:0]   shift_reg_478_re;
  reg        [23:0]   shift_reg_478_im;
  reg        [23:0]   shift_reg_479_re;
  reg        [23:0]   shift_reg_479_im;
  reg        [23:0]   shift_reg_480_re;
  reg        [23:0]   shift_reg_480_im;
  reg        [23:0]   shift_reg_481_re;
  reg        [23:0]   shift_reg_481_im;
  reg        [23:0]   shift_reg_482_re;
  reg        [23:0]   shift_reg_482_im;
  reg        [23:0]   shift_reg_483_re;
  reg        [23:0]   shift_reg_483_im;
  reg        [23:0]   shift_reg_484_re;
  reg        [23:0]   shift_reg_484_im;
  reg        [23:0]   shift_reg_485_re;
  reg        [23:0]   shift_reg_485_im;
  reg        [23:0]   shift_reg_486_re;
  reg        [23:0]   shift_reg_486_im;
  reg        [23:0]   shift_reg_487_re;
  reg        [23:0]   shift_reg_487_im;
  reg        [23:0]   shift_reg_488_re;
  reg        [23:0]   shift_reg_488_im;
  reg        [23:0]   shift_reg_489_re;
  reg        [23:0]   shift_reg_489_im;
  reg        [23:0]   shift_reg_490_re;
  reg        [23:0]   shift_reg_490_im;
  reg        [23:0]   shift_reg_491_re;
  reg        [23:0]   shift_reg_491_im;
  reg        [23:0]   shift_reg_492_re;
  reg        [23:0]   shift_reg_492_im;
  reg        [23:0]   shift_reg_493_re;
  reg        [23:0]   shift_reg_493_im;
  reg        [23:0]   shift_reg_494_re;
  reg        [23:0]   shift_reg_494_im;
  reg        [23:0]   shift_reg_495_re;
  reg        [23:0]   shift_reg_495_im;
  reg        [23:0]   shift_reg_496_re;
  reg        [23:0]   shift_reg_496_im;
  reg        [23:0]   shift_reg_497_re;
  reg        [23:0]   shift_reg_497_im;
  reg        [23:0]   shift_reg_498_re;
  reg        [23:0]   shift_reg_498_im;
  reg        [23:0]   shift_reg_499_re;
  reg        [23:0]   shift_reg_499_im;
  reg        [23:0]   shift_reg_500_re;
  reg        [23:0]   shift_reg_500_im;
  reg        [23:0]   shift_reg_501_re;
  reg        [23:0]   shift_reg_501_im;
  reg        [23:0]   shift_reg_502_re;
  reg        [23:0]   shift_reg_502_im;
  reg        [23:0]   shift_reg_503_re;
  reg        [23:0]   shift_reg_503_im;
  reg        [23:0]   shift_reg_504_re;
  reg        [23:0]   shift_reg_504_im;
  reg        [23:0]   shift_reg_505_re;
  reg        [23:0]   shift_reg_505_im;
  reg        [23:0]   shift_reg_506_re;
  reg        [23:0]   shift_reg_506_im;
  reg        [23:0]   shift_reg_507_re;
  reg        [23:0]   shift_reg_507_im;
  reg        [23:0]   shift_reg_508_re;
  reg        [23:0]   shift_reg_508_im;
  reg        [23:0]   shift_reg_509_re;
  reg        [23:0]   shift_reg_509_im;
  reg        [23:0]   shift_reg_510_re;
  reg        [23:0]   shift_reg_510_im;
  reg        [23:0]   shift_reg_511_re;
  reg        [23:0]   shift_reg_511_im;

  assign output_re = shift_reg_511_re;
  assign output_im = shift_reg_511_im;
  always @(posedge clk) begin
    shift_reg_0_re <= input_re;
    shift_reg_0_im <= input_im;
    shift_reg_1_re <= shift_reg_0_re;
    shift_reg_1_im <= shift_reg_0_im;
    shift_reg_2_re <= shift_reg_1_re;
    shift_reg_2_im <= shift_reg_1_im;
    shift_reg_3_re <= shift_reg_2_re;
    shift_reg_3_im <= shift_reg_2_im;
    shift_reg_4_re <= shift_reg_3_re;
    shift_reg_4_im <= shift_reg_3_im;
    shift_reg_5_re <= shift_reg_4_re;
    shift_reg_5_im <= shift_reg_4_im;
    shift_reg_6_re <= shift_reg_5_re;
    shift_reg_6_im <= shift_reg_5_im;
    shift_reg_7_re <= shift_reg_6_re;
    shift_reg_7_im <= shift_reg_6_im;
    shift_reg_8_re <= shift_reg_7_re;
    shift_reg_8_im <= shift_reg_7_im;
    shift_reg_9_re <= shift_reg_8_re;
    shift_reg_9_im <= shift_reg_8_im;
    shift_reg_10_re <= shift_reg_9_re;
    shift_reg_10_im <= shift_reg_9_im;
    shift_reg_11_re <= shift_reg_10_re;
    shift_reg_11_im <= shift_reg_10_im;
    shift_reg_12_re <= shift_reg_11_re;
    shift_reg_12_im <= shift_reg_11_im;
    shift_reg_13_re <= shift_reg_12_re;
    shift_reg_13_im <= shift_reg_12_im;
    shift_reg_14_re <= shift_reg_13_re;
    shift_reg_14_im <= shift_reg_13_im;
    shift_reg_15_re <= shift_reg_14_re;
    shift_reg_15_im <= shift_reg_14_im;
    shift_reg_16_re <= shift_reg_15_re;
    shift_reg_16_im <= shift_reg_15_im;
    shift_reg_17_re <= shift_reg_16_re;
    shift_reg_17_im <= shift_reg_16_im;
    shift_reg_18_re <= shift_reg_17_re;
    shift_reg_18_im <= shift_reg_17_im;
    shift_reg_19_re <= shift_reg_18_re;
    shift_reg_19_im <= shift_reg_18_im;
    shift_reg_20_re <= shift_reg_19_re;
    shift_reg_20_im <= shift_reg_19_im;
    shift_reg_21_re <= shift_reg_20_re;
    shift_reg_21_im <= shift_reg_20_im;
    shift_reg_22_re <= shift_reg_21_re;
    shift_reg_22_im <= shift_reg_21_im;
    shift_reg_23_re <= shift_reg_22_re;
    shift_reg_23_im <= shift_reg_22_im;
    shift_reg_24_re <= shift_reg_23_re;
    shift_reg_24_im <= shift_reg_23_im;
    shift_reg_25_re <= shift_reg_24_re;
    shift_reg_25_im <= shift_reg_24_im;
    shift_reg_26_re <= shift_reg_25_re;
    shift_reg_26_im <= shift_reg_25_im;
    shift_reg_27_re <= shift_reg_26_re;
    shift_reg_27_im <= shift_reg_26_im;
    shift_reg_28_re <= shift_reg_27_re;
    shift_reg_28_im <= shift_reg_27_im;
    shift_reg_29_re <= shift_reg_28_re;
    shift_reg_29_im <= shift_reg_28_im;
    shift_reg_30_re <= shift_reg_29_re;
    shift_reg_30_im <= shift_reg_29_im;
    shift_reg_31_re <= shift_reg_30_re;
    shift_reg_31_im <= shift_reg_30_im;
    shift_reg_32_re <= shift_reg_31_re;
    shift_reg_32_im <= shift_reg_31_im;
    shift_reg_33_re <= shift_reg_32_re;
    shift_reg_33_im <= shift_reg_32_im;
    shift_reg_34_re <= shift_reg_33_re;
    shift_reg_34_im <= shift_reg_33_im;
    shift_reg_35_re <= shift_reg_34_re;
    shift_reg_35_im <= shift_reg_34_im;
    shift_reg_36_re <= shift_reg_35_re;
    shift_reg_36_im <= shift_reg_35_im;
    shift_reg_37_re <= shift_reg_36_re;
    shift_reg_37_im <= shift_reg_36_im;
    shift_reg_38_re <= shift_reg_37_re;
    shift_reg_38_im <= shift_reg_37_im;
    shift_reg_39_re <= shift_reg_38_re;
    shift_reg_39_im <= shift_reg_38_im;
    shift_reg_40_re <= shift_reg_39_re;
    shift_reg_40_im <= shift_reg_39_im;
    shift_reg_41_re <= shift_reg_40_re;
    shift_reg_41_im <= shift_reg_40_im;
    shift_reg_42_re <= shift_reg_41_re;
    shift_reg_42_im <= shift_reg_41_im;
    shift_reg_43_re <= shift_reg_42_re;
    shift_reg_43_im <= shift_reg_42_im;
    shift_reg_44_re <= shift_reg_43_re;
    shift_reg_44_im <= shift_reg_43_im;
    shift_reg_45_re <= shift_reg_44_re;
    shift_reg_45_im <= shift_reg_44_im;
    shift_reg_46_re <= shift_reg_45_re;
    shift_reg_46_im <= shift_reg_45_im;
    shift_reg_47_re <= shift_reg_46_re;
    shift_reg_47_im <= shift_reg_46_im;
    shift_reg_48_re <= shift_reg_47_re;
    shift_reg_48_im <= shift_reg_47_im;
    shift_reg_49_re <= shift_reg_48_re;
    shift_reg_49_im <= shift_reg_48_im;
    shift_reg_50_re <= shift_reg_49_re;
    shift_reg_50_im <= shift_reg_49_im;
    shift_reg_51_re <= shift_reg_50_re;
    shift_reg_51_im <= shift_reg_50_im;
    shift_reg_52_re <= shift_reg_51_re;
    shift_reg_52_im <= shift_reg_51_im;
    shift_reg_53_re <= shift_reg_52_re;
    shift_reg_53_im <= shift_reg_52_im;
    shift_reg_54_re <= shift_reg_53_re;
    shift_reg_54_im <= shift_reg_53_im;
    shift_reg_55_re <= shift_reg_54_re;
    shift_reg_55_im <= shift_reg_54_im;
    shift_reg_56_re <= shift_reg_55_re;
    shift_reg_56_im <= shift_reg_55_im;
    shift_reg_57_re <= shift_reg_56_re;
    shift_reg_57_im <= shift_reg_56_im;
    shift_reg_58_re <= shift_reg_57_re;
    shift_reg_58_im <= shift_reg_57_im;
    shift_reg_59_re <= shift_reg_58_re;
    shift_reg_59_im <= shift_reg_58_im;
    shift_reg_60_re <= shift_reg_59_re;
    shift_reg_60_im <= shift_reg_59_im;
    shift_reg_61_re <= shift_reg_60_re;
    shift_reg_61_im <= shift_reg_60_im;
    shift_reg_62_re <= shift_reg_61_re;
    shift_reg_62_im <= shift_reg_61_im;
    shift_reg_63_re <= shift_reg_62_re;
    shift_reg_63_im <= shift_reg_62_im;
    shift_reg_64_re <= shift_reg_63_re;
    shift_reg_64_im <= shift_reg_63_im;
    shift_reg_65_re <= shift_reg_64_re;
    shift_reg_65_im <= shift_reg_64_im;
    shift_reg_66_re <= shift_reg_65_re;
    shift_reg_66_im <= shift_reg_65_im;
    shift_reg_67_re <= shift_reg_66_re;
    shift_reg_67_im <= shift_reg_66_im;
    shift_reg_68_re <= shift_reg_67_re;
    shift_reg_68_im <= shift_reg_67_im;
    shift_reg_69_re <= shift_reg_68_re;
    shift_reg_69_im <= shift_reg_68_im;
    shift_reg_70_re <= shift_reg_69_re;
    shift_reg_70_im <= shift_reg_69_im;
    shift_reg_71_re <= shift_reg_70_re;
    shift_reg_71_im <= shift_reg_70_im;
    shift_reg_72_re <= shift_reg_71_re;
    shift_reg_72_im <= shift_reg_71_im;
    shift_reg_73_re <= shift_reg_72_re;
    shift_reg_73_im <= shift_reg_72_im;
    shift_reg_74_re <= shift_reg_73_re;
    shift_reg_74_im <= shift_reg_73_im;
    shift_reg_75_re <= shift_reg_74_re;
    shift_reg_75_im <= shift_reg_74_im;
    shift_reg_76_re <= shift_reg_75_re;
    shift_reg_76_im <= shift_reg_75_im;
    shift_reg_77_re <= shift_reg_76_re;
    shift_reg_77_im <= shift_reg_76_im;
    shift_reg_78_re <= shift_reg_77_re;
    shift_reg_78_im <= shift_reg_77_im;
    shift_reg_79_re <= shift_reg_78_re;
    shift_reg_79_im <= shift_reg_78_im;
    shift_reg_80_re <= shift_reg_79_re;
    shift_reg_80_im <= shift_reg_79_im;
    shift_reg_81_re <= shift_reg_80_re;
    shift_reg_81_im <= shift_reg_80_im;
    shift_reg_82_re <= shift_reg_81_re;
    shift_reg_82_im <= shift_reg_81_im;
    shift_reg_83_re <= shift_reg_82_re;
    shift_reg_83_im <= shift_reg_82_im;
    shift_reg_84_re <= shift_reg_83_re;
    shift_reg_84_im <= shift_reg_83_im;
    shift_reg_85_re <= shift_reg_84_re;
    shift_reg_85_im <= shift_reg_84_im;
    shift_reg_86_re <= shift_reg_85_re;
    shift_reg_86_im <= shift_reg_85_im;
    shift_reg_87_re <= shift_reg_86_re;
    shift_reg_87_im <= shift_reg_86_im;
    shift_reg_88_re <= shift_reg_87_re;
    shift_reg_88_im <= shift_reg_87_im;
    shift_reg_89_re <= shift_reg_88_re;
    shift_reg_89_im <= shift_reg_88_im;
    shift_reg_90_re <= shift_reg_89_re;
    shift_reg_90_im <= shift_reg_89_im;
    shift_reg_91_re <= shift_reg_90_re;
    shift_reg_91_im <= shift_reg_90_im;
    shift_reg_92_re <= shift_reg_91_re;
    shift_reg_92_im <= shift_reg_91_im;
    shift_reg_93_re <= shift_reg_92_re;
    shift_reg_93_im <= shift_reg_92_im;
    shift_reg_94_re <= shift_reg_93_re;
    shift_reg_94_im <= shift_reg_93_im;
    shift_reg_95_re <= shift_reg_94_re;
    shift_reg_95_im <= shift_reg_94_im;
    shift_reg_96_re <= shift_reg_95_re;
    shift_reg_96_im <= shift_reg_95_im;
    shift_reg_97_re <= shift_reg_96_re;
    shift_reg_97_im <= shift_reg_96_im;
    shift_reg_98_re <= shift_reg_97_re;
    shift_reg_98_im <= shift_reg_97_im;
    shift_reg_99_re <= shift_reg_98_re;
    shift_reg_99_im <= shift_reg_98_im;
    shift_reg_100_re <= shift_reg_99_re;
    shift_reg_100_im <= shift_reg_99_im;
    shift_reg_101_re <= shift_reg_100_re;
    shift_reg_101_im <= shift_reg_100_im;
    shift_reg_102_re <= shift_reg_101_re;
    shift_reg_102_im <= shift_reg_101_im;
    shift_reg_103_re <= shift_reg_102_re;
    shift_reg_103_im <= shift_reg_102_im;
    shift_reg_104_re <= shift_reg_103_re;
    shift_reg_104_im <= shift_reg_103_im;
    shift_reg_105_re <= shift_reg_104_re;
    shift_reg_105_im <= shift_reg_104_im;
    shift_reg_106_re <= shift_reg_105_re;
    shift_reg_106_im <= shift_reg_105_im;
    shift_reg_107_re <= shift_reg_106_re;
    shift_reg_107_im <= shift_reg_106_im;
    shift_reg_108_re <= shift_reg_107_re;
    shift_reg_108_im <= shift_reg_107_im;
    shift_reg_109_re <= shift_reg_108_re;
    shift_reg_109_im <= shift_reg_108_im;
    shift_reg_110_re <= shift_reg_109_re;
    shift_reg_110_im <= shift_reg_109_im;
    shift_reg_111_re <= shift_reg_110_re;
    shift_reg_111_im <= shift_reg_110_im;
    shift_reg_112_re <= shift_reg_111_re;
    shift_reg_112_im <= shift_reg_111_im;
    shift_reg_113_re <= shift_reg_112_re;
    shift_reg_113_im <= shift_reg_112_im;
    shift_reg_114_re <= shift_reg_113_re;
    shift_reg_114_im <= shift_reg_113_im;
    shift_reg_115_re <= shift_reg_114_re;
    shift_reg_115_im <= shift_reg_114_im;
    shift_reg_116_re <= shift_reg_115_re;
    shift_reg_116_im <= shift_reg_115_im;
    shift_reg_117_re <= shift_reg_116_re;
    shift_reg_117_im <= shift_reg_116_im;
    shift_reg_118_re <= shift_reg_117_re;
    shift_reg_118_im <= shift_reg_117_im;
    shift_reg_119_re <= shift_reg_118_re;
    shift_reg_119_im <= shift_reg_118_im;
    shift_reg_120_re <= shift_reg_119_re;
    shift_reg_120_im <= shift_reg_119_im;
    shift_reg_121_re <= shift_reg_120_re;
    shift_reg_121_im <= shift_reg_120_im;
    shift_reg_122_re <= shift_reg_121_re;
    shift_reg_122_im <= shift_reg_121_im;
    shift_reg_123_re <= shift_reg_122_re;
    shift_reg_123_im <= shift_reg_122_im;
    shift_reg_124_re <= shift_reg_123_re;
    shift_reg_124_im <= shift_reg_123_im;
    shift_reg_125_re <= shift_reg_124_re;
    shift_reg_125_im <= shift_reg_124_im;
    shift_reg_126_re <= shift_reg_125_re;
    shift_reg_126_im <= shift_reg_125_im;
    shift_reg_127_re <= shift_reg_126_re;
    shift_reg_127_im <= shift_reg_126_im;
    shift_reg_128_re <= shift_reg_127_re;
    shift_reg_128_im <= shift_reg_127_im;
    shift_reg_129_re <= shift_reg_128_re;
    shift_reg_129_im <= shift_reg_128_im;
    shift_reg_130_re <= shift_reg_129_re;
    shift_reg_130_im <= shift_reg_129_im;
    shift_reg_131_re <= shift_reg_130_re;
    shift_reg_131_im <= shift_reg_130_im;
    shift_reg_132_re <= shift_reg_131_re;
    shift_reg_132_im <= shift_reg_131_im;
    shift_reg_133_re <= shift_reg_132_re;
    shift_reg_133_im <= shift_reg_132_im;
    shift_reg_134_re <= shift_reg_133_re;
    shift_reg_134_im <= shift_reg_133_im;
    shift_reg_135_re <= shift_reg_134_re;
    shift_reg_135_im <= shift_reg_134_im;
    shift_reg_136_re <= shift_reg_135_re;
    shift_reg_136_im <= shift_reg_135_im;
    shift_reg_137_re <= shift_reg_136_re;
    shift_reg_137_im <= shift_reg_136_im;
    shift_reg_138_re <= shift_reg_137_re;
    shift_reg_138_im <= shift_reg_137_im;
    shift_reg_139_re <= shift_reg_138_re;
    shift_reg_139_im <= shift_reg_138_im;
    shift_reg_140_re <= shift_reg_139_re;
    shift_reg_140_im <= shift_reg_139_im;
    shift_reg_141_re <= shift_reg_140_re;
    shift_reg_141_im <= shift_reg_140_im;
    shift_reg_142_re <= shift_reg_141_re;
    shift_reg_142_im <= shift_reg_141_im;
    shift_reg_143_re <= shift_reg_142_re;
    shift_reg_143_im <= shift_reg_142_im;
    shift_reg_144_re <= shift_reg_143_re;
    shift_reg_144_im <= shift_reg_143_im;
    shift_reg_145_re <= shift_reg_144_re;
    shift_reg_145_im <= shift_reg_144_im;
    shift_reg_146_re <= shift_reg_145_re;
    shift_reg_146_im <= shift_reg_145_im;
    shift_reg_147_re <= shift_reg_146_re;
    shift_reg_147_im <= shift_reg_146_im;
    shift_reg_148_re <= shift_reg_147_re;
    shift_reg_148_im <= shift_reg_147_im;
    shift_reg_149_re <= shift_reg_148_re;
    shift_reg_149_im <= shift_reg_148_im;
    shift_reg_150_re <= shift_reg_149_re;
    shift_reg_150_im <= shift_reg_149_im;
    shift_reg_151_re <= shift_reg_150_re;
    shift_reg_151_im <= shift_reg_150_im;
    shift_reg_152_re <= shift_reg_151_re;
    shift_reg_152_im <= shift_reg_151_im;
    shift_reg_153_re <= shift_reg_152_re;
    shift_reg_153_im <= shift_reg_152_im;
    shift_reg_154_re <= shift_reg_153_re;
    shift_reg_154_im <= shift_reg_153_im;
    shift_reg_155_re <= shift_reg_154_re;
    shift_reg_155_im <= shift_reg_154_im;
    shift_reg_156_re <= shift_reg_155_re;
    shift_reg_156_im <= shift_reg_155_im;
    shift_reg_157_re <= shift_reg_156_re;
    shift_reg_157_im <= shift_reg_156_im;
    shift_reg_158_re <= shift_reg_157_re;
    shift_reg_158_im <= shift_reg_157_im;
    shift_reg_159_re <= shift_reg_158_re;
    shift_reg_159_im <= shift_reg_158_im;
    shift_reg_160_re <= shift_reg_159_re;
    shift_reg_160_im <= shift_reg_159_im;
    shift_reg_161_re <= shift_reg_160_re;
    shift_reg_161_im <= shift_reg_160_im;
    shift_reg_162_re <= shift_reg_161_re;
    shift_reg_162_im <= shift_reg_161_im;
    shift_reg_163_re <= shift_reg_162_re;
    shift_reg_163_im <= shift_reg_162_im;
    shift_reg_164_re <= shift_reg_163_re;
    shift_reg_164_im <= shift_reg_163_im;
    shift_reg_165_re <= shift_reg_164_re;
    shift_reg_165_im <= shift_reg_164_im;
    shift_reg_166_re <= shift_reg_165_re;
    shift_reg_166_im <= shift_reg_165_im;
    shift_reg_167_re <= shift_reg_166_re;
    shift_reg_167_im <= shift_reg_166_im;
    shift_reg_168_re <= shift_reg_167_re;
    shift_reg_168_im <= shift_reg_167_im;
    shift_reg_169_re <= shift_reg_168_re;
    shift_reg_169_im <= shift_reg_168_im;
    shift_reg_170_re <= shift_reg_169_re;
    shift_reg_170_im <= shift_reg_169_im;
    shift_reg_171_re <= shift_reg_170_re;
    shift_reg_171_im <= shift_reg_170_im;
    shift_reg_172_re <= shift_reg_171_re;
    shift_reg_172_im <= shift_reg_171_im;
    shift_reg_173_re <= shift_reg_172_re;
    shift_reg_173_im <= shift_reg_172_im;
    shift_reg_174_re <= shift_reg_173_re;
    shift_reg_174_im <= shift_reg_173_im;
    shift_reg_175_re <= shift_reg_174_re;
    shift_reg_175_im <= shift_reg_174_im;
    shift_reg_176_re <= shift_reg_175_re;
    shift_reg_176_im <= shift_reg_175_im;
    shift_reg_177_re <= shift_reg_176_re;
    shift_reg_177_im <= shift_reg_176_im;
    shift_reg_178_re <= shift_reg_177_re;
    shift_reg_178_im <= shift_reg_177_im;
    shift_reg_179_re <= shift_reg_178_re;
    shift_reg_179_im <= shift_reg_178_im;
    shift_reg_180_re <= shift_reg_179_re;
    shift_reg_180_im <= shift_reg_179_im;
    shift_reg_181_re <= shift_reg_180_re;
    shift_reg_181_im <= shift_reg_180_im;
    shift_reg_182_re <= shift_reg_181_re;
    shift_reg_182_im <= shift_reg_181_im;
    shift_reg_183_re <= shift_reg_182_re;
    shift_reg_183_im <= shift_reg_182_im;
    shift_reg_184_re <= shift_reg_183_re;
    shift_reg_184_im <= shift_reg_183_im;
    shift_reg_185_re <= shift_reg_184_re;
    shift_reg_185_im <= shift_reg_184_im;
    shift_reg_186_re <= shift_reg_185_re;
    shift_reg_186_im <= shift_reg_185_im;
    shift_reg_187_re <= shift_reg_186_re;
    shift_reg_187_im <= shift_reg_186_im;
    shift_reg_188_re <= shift_reg_187_re;
    shift_reg_188_im <= shift_reg_187_im;
    shift_reg_189_re <= shift_reg_188_re;
    shift_reg_189_im <= shift_reg_188_im;
    shift_reg_190_re <= shift_reg_189_re;
    shift_reg_190_im <= shift_reg_189_im;
    shift_reg_191_re <= shift_reg_190_re;
    shift_reg_191_im <= shift_reg_190_im;
    shift_reg_192_re <= shift_reg_191_re;
    shift_reg_192_im <= shift_reg_191_im;
    shift_reg_193_re <= shift_reg_192_re;
    shift_reg_193_im <= shift_reg_192_im;
    shift_reg_194_re <= shift_reg_193_re;
    shift_reg_194_im <= shift_reg_193_im;
    shift_reg_195_re <= shift_reg_194_re;
    shift_reg_195_im <= shift_reg_194_im;
    shift_reg_196_re <= shift_reg_195_re;
    shift_reg_196_im <= shift_reg_195_im;
    shift_reg_197_re <= shift_reg_196_re;
    shift_reg_197_im <= shift_reg_196_im;
    shift_reg_198_re <= shift_reg_197_re;
    shift_reg_198_im <= shift_reg_197_im;
    shift_reg_199_re <= shift_reg_198_re;
    shift_reg_199_im <= shift_reg_198_im;
    shift_reg_200_re <= shift_reg_199_re;
    shift_reg_200_im <= shift_reg_199_im;
    shift_reg_201_re <= shift_reg_200_re;
    shift_reg_201_im <= shift_reg_200_im;
    shift_reg_202_re <= shift_reg_201_re;
    shift_reg_202_im <= shift_reg_201_im;
    shift_reg_203_re <= shift_reg_202_re;
    shift_reg_203_im <= shift_reg_202_im;
    shift_reg_204_re <= shift_reg_203_re;
    shift_reg_204_im <= shift_reg_203_im;
    shift_reg_205_re <= shift_reg_204_re;
    shift_reg_205_im <= shift_reg_204_im;
    shift_reg_206_re <= shift_reg_205_re;
    shift_reg_206_im <= shift_reg_205_im;
    shift_reg_207_re <= shift_reg_206_re;
    shift_reg_207_im <= shift_reg_206_im;
    shift_reg_208_re <= shift_reg_207_re;
    shift_reg_208_im <= shift_reg_207_im;
    shift_reg_209_re <= shift_reg_208_re;
    shift_reg_209_im <= shift_reg_208_im;
    shift_reg_210_re <= shift_reg_209_re;
    shift_reg_210_im <= shift_reg_209_im;
    shift_reg_211_re <= shift_reg_210_re;
    shift_reg_211_im <= shift_reg_210_im;
    shift_reg_212_re <= shift_reg_211_re;
    shift_reg_212_im <= shift_reg_211_im;
    shift_reg_213_re <= shift_reg_212_re;
    shift_reg_213_im <= shift_reg_212_im;
    shift_reg_214_re <= shift_reg_213_re;
    shift_reg_214_im <= shift_reg_213_im;
    shift_reg_215_re <= shift_reg_214_re;
    shift_reg_215_im <= shift_reg_214_im;
    shift_reg_216_re <= shift_reg_215_re;
    shift_reg_216_im <= shift_reg_215_im;
    shift_reg_217_re <= shift_reg_216_re;
    shift_reg_217_im <= shift_reg_216_im;
    shift_reg_218_re <= shift_reg_217_re;
    shift_reg_218_im <= shift_reg_217_im;
    shift_reg_219_re <= shift_reg_218_re;
    shift_reg_219_im <= shift_reg_218_im;
    shift_reg_220_re <= shift_reg_219_re;
    shift_reg_220_im <= shift_reg_219_im;
    shift_reg_221_re <= shift_reg_220_re;
    shift_reg_221_im <= shift_reg_220_im;
    shift_reg_222_re <= shift_reg_221_re;
    shift_reg_222_im <= shift_reg_221_im;
    shift_reg_223_re <= shift_reg_222_re;
    shift_reg_223_im <= shift_reg_222_im;
    shift_reg_224_re <= shift_reg_223_re;
    shift_reg_224_im <= shift_reg_223_im;
    shift_reg_225_re <= shift_reg_224_re;
    shift_reg_225_im <= shift_reg_224_im;
    shift_reg_226_re <= shift_reg_225_re;
    shift_reg_226_im <= shift_reg_225_im;
    shift_reg_227_re <= shift_reg_226_re;
    shift_reg_227_im <= shift_reg_226_im;
    shift_reg_228_re <= shift_reg_227_re;
    shift_reg_228_im <= shift_reg_227_im;
    shift_reg_229_re <= shift_reg_228_re;
    shift_reg_229_im <= shift_reg_228_im;
    shift_reg_230_re <= shift_reg_229_re;
    shift_reg_230_im <= shift_reg_229_im;
    shift_reg_231_re <= shift_reg_230_re;
    shift_reg_231_im <= shift_reg_230_im;
    shift_reg_232_re <= shift_reg_231_re;
    shift_reg_232_im <= shift_reg_231_im;
    shift_reg_233_re <= shift_reg_232_re;
    shift_reg_233_im <= shift_reg_232_im;
    shift_reg_234_re <= shift_reg_233_re;
    shift_reg_234_im <= shift_reg_233_im;
    shift_reg_235_re <= shift_reg_234_re;
    shift_reg_235_im <= shift_reg_234_im;
    shift_reg_236_re <= shift_reg_235_re;
    shift_reg_236_im <= shift_reg_235_im;
    shift_reg_237_re <= shift_reg_236_re;
    shift_reg_237_im <= shift_reg_236_im;
    shift_reg_238_re <= shift_reg_237_re;
    shift_reg_238_im <= shift_reg_237_im;
    shift_reg_239_re <= shift_reg_238_re;
    shift_reg_239_im <= shift_reg_238_im;
    shift_reg_240_re <= shift_reg_239_re;
    shift_reg_240_im <= shift_reg_239_im;
    shift_reg_241_re <= shift_reg_240_re;
    shift_reg_241_im <= shift_reg_240_im;
    shift_reg_242_re <= shift_reg_241_re;
    shift_reg_242_im <= shift_reg_241_im;
    shift_reg_243_re <= shift_reg_242_re;
    shift_reg_243_im <= shift_reg_242_im;
    shift_reg_244_re <= shift_reg_243_re;
    shift_reg_244_im <= shift_reg_243_im;
    shift_reg_245_re <= shift_reg_244_re;
    shift_reg_245_im <= shift_reg_244_im;
    shift_reg_246_re <= shift_reg_245_re;
    shift_reg_246_im <= shift_reg_245_im;
    shift_reg_247_re <= shift_reg_246_re;
    shift_reg_247_im <= shift_reg_246_im;
    shift_reg_248_re <= shift_reg_247_re;
    shift_reg_248_im <= shift_reg_247_im;
    shift_reg_249_re <= shift_reg_248_re;
    shift_reg_249_im <= shift_reg_248_im;
    shift_reg_250_re <= shift_reg_249_re;
    shift_reg_250_im <= shift_reg_249_im;
    shift_reg_251_re <= shift_reg_250_re;
    shift_reg_251_im <= shift_reg_250_im;
    shift_reg_252_re <= shift_reg_251_re;
    shift_reg_252_im <= shift_reg_251_im;
    shift_reg_253_re <= shift_reg_252_re;
    shift_reg_253_im <= shift_reg_252_im;
    shift_reg_254_re <= shift_reg_253_re;
    shift_reg_254_im <= shift_reg_253_im;
    shift_reg_255_re <= shift_reg_254_re;
    shift_reg_255_im <= shift_reg_254_im;
    shift_reg_256_re <= shift_reg_255_re;
    shift_reg_256_im <= shift_reg_255_im;
    shift_reg_257_re <= shift_reg_256_re;
    shift_reg_257_im <= shift_reg_256_im;
    shift_reg_258_re <= shift_reg_257_re;
    shift_reg_258_im <= shift_reg_257_im;
    shift_reg_259_re <= shift_reg_258_re;
    shift_reg_259_im <= shift_reg_258_im;
    shift_reg_260_re <= shift_reg_259_re;
    shift_reg_260_im <= shift_reg_259_im;
    shift_reg_261_re <= shift_reg_260_re;
    shift_reg_261_im <= shift_reg_260_im;
    shift_reg_262_re <= shift_reg_261_re;
    shift_reg_262_im <= shift_reg_261_im;
    shift_reg_263_re <= shift_reg_262_re;
    shift_reg_263_im <= shift_reg_262_im;
    shift_reg_264_re <= shift_reg_263_re;
    shift_reg_264_im <= shift_reg_263_im;
    shift_reg_265_re <= shift_reg_264_re;
    shift_reg_265_im <= shift_reg_264_im;
    shift_reg_266_re <= shift_reg_265_re;
    shift_reg_266_im <= shift_reg_265_im;
    shift_reg_267_re <= shift_reg_266_re;
    shift_reg_267_im <= shift_reg_266_im;
    shift_reg_268_re <= shift_reg_267_re;
    shift_reg_268_im <= shift_reg_267_im;
    shift_reg_269_re <= shift_reg_268_re;
    shift_reg_269_im <= shift_reg_268_im;
    shift_reg_270_re <= shift_reg_269_re;
    shift_reg_270_im <= shift_reg_269_im;
    shift_reg_271_re <= shift_reg_270_re;
    shift_reg_271_im <= shift_reg_270_im;
    shift_reg_272_re <= shift_reg_271_re;
    shift_reg_272_im <= shift_reg_271_im;
    shift_reg_273_re <= shift_reg_272_re;
    shift_reg_273_im <= shift_reg_272_im;
    shift_reg_274_re <= shift_reg_273_re;
    shift_reg_274_im <= shift_reg_273_im;
    shift_reg_275_re <= shift_reg_274_re;
    shift_reg_275_im <= shift_reg_274_im;
    shift_reg_276_re <= shift_reg_275_re;
    shift_reg_276_im <= shift_reg_275_im;
    shift_reg_277_re <= shift_reg_276_re;
    shift_reg_277_im <= shift_reg_276_im;
    shift_reg_278_re <= shift_reg_277_re;
    shift_reg_278_im <= shift_reg_277_im;
    shift_reg_279_re <= shift_reg_278_re;
    shift_reg_279_im <= shift_reg_278_im;
    shift_reg_280_re <= shift_reg_279_re;
    shift_reg_280_im <= shift_reg_279_im;
    shift_reg_281_re <= shift_reg_280_re;
    shift_reg_281_im <= shift_reg_280_im;
    shift_reg_282_re <= shift_reg_281_re;
    shift_reg_282_im <= shift_reg_281_im;
    shift_reg_283_re <= shift_reg_282_re;
    shift_reg_283_im <= shift_reg_282_im;
    shift_reg_284_re <= shift_reg_283_re;
    shift_reg_284_im <= shift_reg_283_im;
    shift_reg_285_re <= shift_reg_284_re;
    shift_reg_285_im <= shift_reg_284_im;
    shift_reg_286_re <= shift_reg_285_re;
    shift_reg_286_im <= shift_reg_285_im;
    shift_reg_287_re <= shift_reg_286_re;
    shift_reg_287_im <= shift_reg_286_im;
    shift_reg_288_re <= shift_reg_287_re;
    shift_reg_288_im <= shift_reg_287_im;
    shift_reg_289_re <= shift_reg_288_re;
    shift_reg_289_im <= shift_reg_288_im;
    shift_reg_290_re <= shift_reg_289_re;
    shift_reg_290_im <= shift_reg_289_im;
    shift_reg_291_re <= shift_reg_290_re;
    shift_reg_291_im <= shift_reg_290_im;
    shift_reg_292_re <= shift_reg_291_re;
    shift_reg_292_im <= shift_reg_291_im;
    shift_reg_293_re <= shift_reg_292_re;
    shift_reg_293_im <= shift_reg_292_im;
    shift_reg_294_re <= shift_reg_293_re;
    shift_reg_294_im <= shift_reg_293_im;
    shift_reg_295_re <= shift_reg_294_re;
    shift_reg_295_im <= shift_reg_294_im;
    shift_reg_296_re <= shift_reg_295_re;
    shift_reg_296_im <= shift_reg_295_im;
    shift_reg_297_re <= shift_reg_296_re;
    shift_reg_297_im <= shift_reg_296_im;
    shift_reg_298_re <= shift_reg_297_re;
    shift_reg_298_im <= shift_reg_297_im;
    shift_reg_299_re <= shift_reg_298_re;
    shift_reg_299_im <= shift_reg_298_im;
    shift_reg_300_re <= shift_reg_299_re;
    shift_reg_300_im <= shift_reg_299_im;
    shift_reg_301_re <= shift_reg_300_re;
    shift_reg_301_im <= shift_reg_300_im;
    shift_reg_302_re <= shift_reg_301_re;
    shift_reg_302_im <= shift_reg_301_im;
    shift_reg_303_re <= shift_reg_302_re;
    shift_reg_303_im <= shift_reg_302_im;
    shift_reg_304_re <= shift_reg_303_re;
    shift_reg_304_im <= shift_reg_303_im;
    shift_reg_305_re <= shift_reg_304_re;
    shift_reg_305_im <= shift_reg_304_im;
    shift_reg_306_re <= shift_reg_305_re;
    shift_reg_306_im <= shift_reg_305_im;
    shift_reg_307_re <= shift_reg_306_re;
    shift_reg_307_im <= shift_reg_306_im;
    shift_reg_308_re <= shift_reg_307_re;
    shift_reg_308_im <= shift_reg_307_im;
    shift_reg_309_re <= shift_reg_308_re;
    shift_reg_309_im <= shift_reg_308_im;
    shift_reg_310_re <= shift_reg_309_re;
    shift_reg_310_im <= shift_reg_309_im;
    shift_reg_311_re <= shift_reg_310_re;
    shift_reg_311_im <= shift_reg_310_im;
    shift_reg_312_re <= shift_reg_311_re;
    shift_reg_312_im <= shift_reg_311_im;
    shift_reg_313_re <= shift_reg_312_re;
    shift_reg_313_im <= shift_reg_312_im;
    shift_reg_314_re <= shift_reg_313_re;
    shift_reg_314_im <= shift_reg_313_im;
    shift_reg_315_re <= shift_reg_314_re;
    shift_reg_315_im <= shift_reg_314_im;
    shift_reg_316_re <= shift_reg_315_re;
    shift_reg_316_im <= shift_reg_315_im;
    shift_reg_317_re <= shift_reg_316_re;
    shift_reg_317_im <= shift_reg_316_im;
    shift_reg_318_re <= shift_reg_317_re;
    shift_reg_318_im <= shift_reg_317_im;
    shift_reg_319_re <= shift_reg_318_re;
    shift_reg_319_im <= shift_reg_318_im;
    shift_reg_320_re <= shift_reg_319_re;
    shift_reg_320_im <= shift_reg_319_im;
    shift_reg_321_re <= shift_reg_320_re;
    shift_reg_321_im <= shift_reg_320_im;
    shift_reg_322_re <= shift_reg_321_re;
    shift_reg_322_im <= shift_reg_321_im;
    shift_reg_323_re <= shift_reg_322_re;
    shift_reg_323_im <= shift_reg_322_im;
    shift_reg_324_re <= shift_reg_323_re;
    shift_reg_324_im <= shift_reg_323_im;
    shift_reg_325_re <= shift_reg_324_re;
    shift_reg_325_im <= shift_reg_324_im;
    shift_reg_326_re <= shift_reg_325_re;
    shift_reg_326_im <= shift_reg_325_im;
    shift_reg_327_re <= shift_reg_326_re;
    shift_reg_327_im <= shift_reg_326_im;
    shift_reg_328_re <= shift_reg_327_re;
    shift_reg_328_im <= shift_reg_327_im;
    shift_reg_329_re <= shift_reg_328_re;
    shift_reg_329_im <= shift_reg_328_im;
    shift_reg_330_re <= shift_reg_329_re;
    shift_reg_330_im <= shift_reg_329_im;
    shift_reg_331_re <= shift_reg_330_re;
    shift_reg_331_im <= shift_reg_330_im;
    shift_reg_332_re <= shift_reg_331_re;
    shift_reg_332_im <= shift_reg_331_im;
    shift_reg_333_re <= shift_reg_332_re;
    shift_reg_333_im <= shift_reg_332_im;
    shift_reg_334_re <= shift_reg_333_re;
    shift_reg_334_im <= shift_reg_333_im;
    shift_reg_335_re <= shift_reg_334_re;
    shift_reg_335_im <= shift_reg_334_im;
    shift_reg_336_re <= shift_reg_335_re;
    shift_reg_336_im <= shift_reg_335_im;
    shift_reg_337_re <= shift_reg_336_re;
    shift_reg_337_im <= shift_reg_336_im;
    shift_reg_338_re <= shift_reg_337_re;
    shift_reg_338_im <= shift_reg_337_im;
    shift_reg_339_re <= shift_reg_338_re;
    shift_reg_339_im <= shift_reg_338_im;
    shift_reg_340_re <= shift_reg_339_re;
    shift_reg_340_im <= shift_reg_339_im;
    shift_reg_341_re <= shift_reg_340_re;
    shift_reg_341_im <= shift_reg_340_im;
    shift_reg_342_re <= shift_reg_341_re;
    shift_reg_342_im <= shift_reg_341_im;
    shift_reg_343_re <= shift_reg_342_re;
    shift_reg_343_im <= shift_reg_342_im;
    shift_reg_344_re <= shift_reg_343_re;
    shift_reg_344_im <= shift_reg_343_im;
    shift_reg_345_re <= shift_reg_344_re;
    shift_reg_345_im <= shift_reg_344_im;
    shift_reg_346_re <= shift_reg_345_re;
    shift_reg_346_im <= shift_reg_345_im;
    shift_reg_347_re <= shift_reg_346_re;
    shift_reg_347_im <= shift_reg_346_im;
    shift_reg_348_re <= shift_reg_347_re;
    shift_reg_348_im <= shift_reg_347_im;
    shift_reg_349_re <= shift_reg_348_re;
    shift_reg_349_im <= shift_reg_348_im;
    shift_reg_350_re <= shift_reg_349_re;
    shift_reg_350_im <= shift_reg_349_im;
    shift_reg_351_re <= shift_reg_350_re;
    shift_reg_351_im <= shift_reg_350_im;
    shift_reg_352_re <= shift_reg_351_re;
    shift_reg_352_im <= shift_reg_351_im;
    shift_reg_353_re <= shift_reg_352_re;
    shift_reg_353_im <= shift_reg_352_im;
    shift_reg_354_re <= shift_reg_353_re;
    shift_reg_354_im <= shift_reg_353_im;
    shift_reg_355_re <= shift_reg_354_re;
    shift_reg_355_im <= shift_reg_354_im;
    shift_reg_356_re <= shift_reg_355_re;
    shift_reg_356_im <= shift_reg_355_im;
    shift_reg_357_re <= shift_reg_356_re;
    shift_reg_357_im <= shift_reg_356_im;
    shift_reg_358_re <= shift_reg_357_re;
    shift_reg_358_im <= shift_reg_357_im;
    shift_reg_359_re <= shift_reg_358_re;
    shift_reg_359_im <= shift_reg_358_im;
    shift_reg_360_re <= shift_reg_359_re;
    shift_reg_360_im <= shift_reg_359_im;
    shift_reg_361_re <= shift_reg_360_re;
    shift_reg_361_im <= shift_reg_360_im;
    shift_reg_362_re <= shift_reg_361_re;
    shift_reg_362_im <= shift_reg_361_im;
    shift_reg_363_re <= shift_reg_362_re;
    shift_reg_363_im <= shift_reg_362_im;
    shift_reg_364_re <= shift_reg_363_re;
    shift_reg_364_im <= shift_reg_363_im;
    shift_reg_365_re <= shift_reg_364_re;
    shift_reg_365_im <= shift_reg_364_im;
    shift_reg_366_re <= shift_reg_365_re;
    shift_reg_366_im <= shift_reg_365_im;
    shift_reg_367_re <= shift_reg_366_re;
    shift_reg_367_im <= shift_reg_366_im;
    shift_reg_368_re <= shift_reg_367_re;
    shift_reg_368_im <= shift_reg_367_im;
    shift_reg_369_re <= shift_reg_368_re;
    shift_reg_369_im <= shift_reg_368_im;
    shift_reg_370_re <= shift_reg_369_re;
    shift_reg_370_im <= shift_reg_369_im;
    shift_reg_371_re <= shift_reg_370_re;
    shift_reg_371_im <= shift_reg_370_im;
    shift_reg_372_re <= shift_reg_371_re;
    shift_reg_372_im <= shift_reg_371_im;
    shift_reg_373_re <= shift_reg_372_re;
    shift_reg_373_im <= shift_reg_372_im;
    shift_reg_374_re <= shift_reg_373_re;
    shift_reg_374_im <= shift_reg_373_im;
    shift_reg_375_re <= shift_reg_374_re;
    shift_reg_375_im <= shift_reg_374_im;
    shift_reg_376_re <= shift_reg_375_re;
    shift_reg_376_im <= shift_reg_375_im;
    shift_reg_377_re <= shift_reg_376_re;
    shift_reg_377_im <= shift_reg_376_im;
    shift_reg_378_re <= shift_reg_377_re;
    shift_reg_378_im <= shift_reg_377_im;
    shift_reg_379_re <= shift_reg_378_re;
    shift_reg_379_im <= shift_reg_378_im;
    shift_reg_380_re <= shift_reg_379_re;
    shift_reg_380_im <= shift_reg_379_im;
    shift_reg_381_re <= shift_reg_380_re;
    shift_reg_381_im <= shift_reg_380_im;
    shift_reg_382_re <= shift_reg_381_re;
    shift_reg_382_im <= shift_reg_381_im;
    shift_reg_383_re <= shift_reg_382_re;
    shift_reg_383_im <= shift_reg_382_im;
    shift_reg_384_re <= shift_reg_383_re;
    shift_reg_384_im <= shift_reg_383_im;
    shift_reg_385_re <= shift_reg_384_re;
    shift_reg_385_im <= shift_reg_384_im;
    shift_reg_386_re <= shift_reg_385_re;
    shift_reg_386_im <= shift_reg_385_im;
    shift_reg_387_re <= shift_reg_386_re;
    shift_reg_387_im <= shift_reg_386_im;
    shift_reg_388_re <= shift_reg_387_re;
    shift_reg_388_im <= shift_reg_387_im;
    shift_reg_389_re <= shift_reg_388_re;
    shift_reg_389_im <= shift_reg_388_im;
    shift_reg_390_re <= shift_reg_389_re;
    shift_reg_390_im <= shift_reg_389_im;
    shift_reg_391_re <= shift_reg_390_re;
    shift_reg_391_im <= shift_reg_390_im;
    shift_reg_392_re <= shift_reg_391_re;
    shift_reg_392_im <= shift_reg_391_im;
    shift_reg_393_re <= shift_reg_392_re;
    shift_reg_393_im <= shift_reg_392_im;
    shift_reg_394_re <= shift_reg_393_re;
    shift_reg_394_im <= shift_reg_393_im;
    shift_reg_395_re <= shift_reg_394_re;
    shift_reg_395_im <= shift_reg_394_im;
    shift_reg_396_re <= shift_reg_395_re;
    shift_reg_396_im <= shift_reg_395_im;
    shift_reg_397_re <= shift_reg_396_re;
    shift_reg_397_im <= shift_reg_396_im;
    shift_reg_398_re <= shift_reg_397_re;
    shift_reg_398_im <= shift_reg_397_im;
    shift_reg_399_re <= shift_reg_398_re;
    shift_reg_399_im <= shift_reg_398_im;
    shift_reg_400_re <= shift_reg_399_re;
    shift_reg_400_im <= shift_reg_399_im;
    shift_reg_401_re <= shift_reg_400_re;
    shift_reg_401_im <= shift_reg_400_im;
    shift_reg_402_re <= shift_reg_401_re;
    shift_reg_402_im <= shift_reg_401_im;
    shift_reg_403_re <= shift_reg_402_re;
    shift_reg_403_im <= shift_reg_402_im;
    shift_reg_404_re <= shift_reg_403_re;
    shift_reg_404_im <= shift_reg_403_im;
    shift_reg_405_re <= shift_reg_404_re;
    shift_reg_405_im <= shift_reg_404_im;
    shift_reg_406_re <= shift_reg_405_re;
    shift_reg_406_im <= shift_reg_405_im;
    shift_reg_407_re <= shift_reg_406_re;
    shift_reg_407_im <= shift_reg_406_im;
    shift_reg_408_re <= shift_reg_407_re;
    shift_reg_408_im <= shift_reg_407_im;
    shift_reg_409_re <= shift_reg_408_re;
    shift_reg_409_im <= shift_reg_408_im;
    shift_reg_410_re <= shift_reg_409_re;
    shift_reg_410_im <= shift_reg_409_im;
    shift_reg_411_re <= shift_reg_410_re;
    shift_reg_411_im <= shift_reg_410_im;
    shift_reg_412_re <= shift_reg_411_re;
    shift_reg_412_im <= shift_reg_411_im;
    shift_reg_413_re <= shift_reg_412_re;
    shift_reg_413_im <= shift_reg_412_im;
    shift_reg_414_re <= shift_reg_413_re;
    shift_reg_414_im <= shift_reg_413_im;
    shift_reg_415_re <= shift_reg_414_re;
    shift_reg_415_im <= shift_reg_414_im;
    shift_reg_416_re <= shift_reg_415_re;
    shift_reg_416_im <= shift_reg_415_im;
    shift_reg_417_re <= shift_reg_416_re;
    shift_reg_417_im <= shift_reg_416_im;
    shift_reg_418_re <= shift_reg_417_re;
    shift_reg_418_im <= shift_reg_417_im;
    shift_reg_419_re <= shift_reg_418_re;
    shift_reg_419_im <= shift_reg_418_im;
    shift_reg_420_re <= shift_reg_419_re;
    shift_reg_420_im <= shift_reg_419_im;
    shift_reg_421_re <= shift_reg_420_re;
    shift_reg_421_im <= shift_reg_420_im;
    shift_reg_422_re <= shift_reg_421_re;
    shift_reg_422_im <= shift_reg_421_im;
    shift_reg_423_re <= shift_reg_422_re;
    shift_reg_423_im <= shift_reg_422_im;
    shift_reg_424_re <= shift_reg_423_re;
    shift_reg_424_im <= shift_reg_423_im;
    shift_reg_425_re <= shift_reg_424_re;
    shift_reg_425_im <= shift_reg_424_im;
    shift_reg_426_re <= shift_reg_425_re;
    shift_reg_426_im <= shift_reg_425_im;
    shift_reg_427_re <= shift_reg_426_re;
    shift_reg_427_im <= shift_reg_426_im;
    shift_reg_428_re <= shift_reg_427_re;
    shift_reg_428_im <= shift_reg_427_im;
    shift_reg_429_re <= shift_reg_428_re;
    shift_reg_429_im <= shift_reg_428_im;
    shift_reg_430_re <= shift_reg_429_re;
    shift_reg_430_im <= shift_reg_429_im;
    shift_reg_431_re <= shift_reg_430_re;
    shift_reg_431_im <= shift_reg_430_im;
    shift_reg_432_re <= shift_reg_431_re;
    shift_reg_432_im <= shift_reg_431_im;
    shift_reg_433_re <= shift_reg_432_re;
    shift_reg_433_im <= shift_reg_432_im;
    shift_reg_434_re <= shift_reg_433_re;
    shift_reg_434_im <= shift_reg_433_im;
    shift_reg_435_re <= shift_reg_434_re;
    shift_reg_435_im <= shift_reg_434_im;
    shift_reg_436_re <= shift_reg_435_re;
    shift_reg_436_im <= shift_reg_435_im;
    shift_reg_437_re <= shift_reg_436_re;
    shift_reg_437_im <= shift_reg_436_im;
    shift_reg_438_re <= shift_reg_437_re;
    shift_reg_438_im <= shift_reg_437_im;
    shift_reg_439_re <= shift_reg_438_re;
    shift_reg_439_im <= shift_reg_438_im;
    shift_reg_440_re <= shift_reg_439_re;
    shift_reg_440_im <= shift_reg_439_im;
    shift_reg_441_re <= shift_reg_440_re;
    shift_reg_441_im <= shift_reg_440_im;
    shift_reg_442_re <= shift_reg_441_re;
    shift_reg_442_im <= shift_reg_441_im;
    shift_reg_443_re <= shift_reg_442_re;
    shift_reg_443_im <= shift_reg_442_im;
    shift_reg_444_re <= shift_reg_443_re;
    shift_reg_444_im <= shift_reg_443_im;
    shift_reg_445_re <= shift_reg_444_re;
    shift_reg_445_im <= shift_reg_444_im;
    shift_reg_446_re <= shift_reg_445_re;
    shift_reg_446_im <= shift_reg_445_im;
    shift_reg_447_re <= shift_reg_446_re;
    shift_reg_447_im <= shift_reg_446_im;
    shift_reg_448_re <= shift_reg_447_re;
    shift_reg_448_im <= shift_reg_447_im;
    shift_reg_449_re <= shift_reg_448_re;
    shift_reg_449_im <= shift_reg_448_im;
    shift_reg_450_re <= shift_reg_449_re;
    shift_reg_450_im <= shift_reg_449_im;
    shift_reg_451_re <= shift_reg_450_re;
    shift_reg_451_im <= shift_reg_450_im;
    shift_reg_452_re <= shift_reg_451_re;
    shift_reg_452_im <= shift_reg_451_im;
    shift_reg_453_re <= shift_reg_452_re;
    shift_reg_453_im <= shift_reg_452_im;
    shift_reg_454_re <= shift_reg_453_re;
    shift_reg_454_im <= shift_reg_453_im;
    shift_reg_455_re <= shift_reg_454_re;
    shift_reg_455_im <= shift_reg_454_im;
    shift_reg_456_re <= shift_reg_455_re;
    shift_reg_456_im <= shift_reg_455_im;
    shift_reg_457_re <= shift_reg_456_re;
    shift_reg_457_im <= shift_reg_456_im;
    shift_reg_458_re <= shift_reg_457_re;
    shift_reg_458_im <= shift_reg_457_im;
    shift_reg_459_re <= shift_reg_458_re;
    shift_reg_459_im <= shift_reg_458_im;
    shift_reg_460_re <= shift_reg_459_re;
    shift_reg_460_im <= shift_reg_459_im;
    shift_reg_461_re <= shift_reg_460_re;
    shift_reg_461_im <= shift_reg_460_im;
    shift_reg_462_re <= shift_reg_461_re;
    shift_reg_462_im <= shift_reg_461_im;
    shift_reg_463_re <= shift_reg_462_re;
    shift_reg_463_im <= shift_reg_462_im;
    shift_reg_464_re <= shift_reg_463_re;
    shift_reg_464_im <= shift_reg_463_im;
    shift_reg_465_re <= shift_reg_464_re;
    shift_reg_465_im <= shift_reg_464_im;
    shift_reg_466_re <= shift_reg_465_re;
    shift_reg_466_im <= shift_reg_465_im;
    shift_reg_467_re <= shift_reg_466_re;
    shift_reg_467_im <= shift_reg_466_im;
    shift_reg_468_re <= shift_reg_467_re;
    shift_reg_468_im <= shift_reg_467_im;
    shift_reg_469_re <= shift_reg_468_re;
    shift_reg_469_im <= shift_reg_468_im;
    shift_reg_470_re <= shift_reg_469_re;
    shift_reg_470_im <= shift_reg_469_im;
    shift_reg_471_re <= shift_reg_470_re;
    shift_reg_471_im <= shift_reg_470_im;
    shift_reg_472_re <= shift_reg_471_re;
    shift_reg_472_im <= shift_reg_471_im;
    shift_reg_473_re <= shift_reg_472_re;
    shift_reg_473_im <= shift_reg_472_im;
    shift_reg_474_re <= shift_reg_473_re;
    shift_reg_474_im <= shift_reg_473_im;
    shift_reg_475_re <= shift_reg_474_re;
    shift_reg_475_im <= shift_reg_474_im;
    shift_reg_476_re <= shift_reg_475_re;
    shift_reg_476_im <= shift_reg_475_im;
    shift_reg_477_re <= shift_reg_476_re;
    shift_reg_477_im <= shift_reg_476_im;
    shift_reg_478_re <= shift_reg_477_re;
    shift_reg_478_im <= shift_reg_477_im;
    shift_reg_479_re <= shift_reg_478_re;
    shift_reg_479_im <= shift_reg_478_im;
    shift_reg_480_re <= shift_reg_479_re;
    shift_reg_480_im <= shift_reg_479_im;
    shift_reg_481_re <= shift_reg_480_re;
    shift_reg_481_im <= shift_reg_480_im;
    shift_reg_482_re <= shift_reg_481_re;
    shift_reg_482_im <= shift_reg_481_im;
    shift_reg_483_re <= shift_reg_482_re;
    shift_reg_483_im <= shift_reg_482_im;
    shift_reg_484_re <= shift_reg_483_re;
    shift_reg_484_im <= shift_reg_483_im;
    shift_reg_485_re <= shift_reg_484_re;
    shift_reg_485_im <= shift_reg_484_im;
    shift_reg_486_re <= shift_reg_485_re;
    shift_reg_486_im <= shift_reg_485_im;
    shift_reg_487_re <= shift_reg_486_re;
    shift_reg_487_im <= shift_reg_486_im;
    shift_reg_488_re <= shift_reg_487_re;
    shift_reg_488_im <= shift_reg_487_im;
    shift_reg_489_re <= shift_reg_488_re;
    shift_reg_489_im <= shift_reg_488_im;
    shift_reg_490_re <= shift_reg_489_re;
    shift_reg_490_im <= shift_reg_489_im;
    shift_reg_491_re <= shift_reg_490_re;
    shift_reg_491_im <= shift_reg_490_im;
    shift_reg_492_re <= shift_reg_491_re;
    shift_reg_492_im <= shift_reg_491_im;
    shift_reg_493_re <= shift_reg_492_re;
    shift_reg_493_im <= shift_reg_492_im;
    shift_reg_494_re <= shift_reg_493_re;
    shift_reg_494_im <= shift_reg_493_im;
    shift_reg_495_re <= shift_reg_494_re;
    shift_reg_495_im <= shift_reg_494_im;
    shift_reg_496_re <= shift_reg_495_re;
    shift_reg_496_im <= shift_reg_495_im;
    shift_reg_497_re <= shift_reg_496_re;
    shift_reg_497_im <= shift_reg_496_im;
    shift_reg_498_re <= shift_reg_497_re;
    shift_reg_498_im <= shift_reg_497_im;
    shift_reg_499_re <= shift_reg_498_re;
    shift_reg_499_im <= shift_reg_498_im;
    shift_reg_500_re <= shift_reg_499_re;
    shift_reg_500_im <= shift_reg_499_im;
    shift_reg_501_re <= shift_reg_500_re;
    shift_reg_501_im <= shift_reg_500_im;
    shift_reg_502_re <= shift_reg_501_re;
    shift_reg_502_im <= shift_reg_501_im;
    shift_reg_503_re <= shift_reg_502_re;
    shift_reg_503_im <= shift_reg_502_im;
    shift_reg_504_re <= shift_reg_503_re;
    shift_reg_504_im <= shift_reg_503_im;
    shift_reg_505_re <= shift_reg_504_re;
    shift_reg_505_im <= shift_reg_504_im;
    shift_reg_506_re <= shift_reg_505_re;
    shift_reg_506_im <= shift_reg_505_im;
    shift_reg_507_re <= shift_reg_506_re;
    shift_reg_507_im <= shift_reg_506_im;
    shift_reg_508_re <= shift_reg_507_re;
    shift_reg_508_im <= shift_reg_507_im;
    shift_reg_509_re <= shift_reg_508_re;
    shift_reg_509_im <= shift_reg_508_im;
    shift_reg_510_re <= shift_reg_509_re;
    shift_reg_510_im <= shift_reg_509_im;
    shift_reg_511_re <= shift_reg_510_re;
    shift_reg_511_im <= shift_reg_510_im;
  end


endmodule

module R2Butterfly (
  input      [23:0]   in1_re,
  input      [23:0]   in1_im,
  input      [23:0]   in2_re,
  input      [23:0]   in2_im,
  input      [23:0]   wn_re,
  input      [23:0]   wn_im,
  output     [23:0]   out1_re,
  output     [23:0]   out1_im,
  output     [23:0]   out2_re,
  output     [23:0]   out2_im
);
  wire       [36:0]   _zz_mul_result_re;
  wire       [47:0]   _zz_mul_result_re_1;
  wire       [47:0]   _zz_mul_result_re_2;
  wire       [47:0]   _zz_mul_result_re_3;
  wire       [36:0]   _zz_mul_result_im;
  wire       [47:0]   _zz_mul_result_im_1;
  wire       [47:0]   _zz_mul_result_im_2;
  wire       [47:0]   _zz_mul_result_im_3;
  wire       [23:0]   add_result_re;
  wire       [23:0]   add_result_im;
  wire       [23:0]   sub_result_re;
  wire       [23:0]   sub_result_im;
  wire       [23:0]   mul_result_re;
  wire       [23:0]   mul_result_im;

  assign _zz_mul_result_re = (_zz_mul_result_re_1 >>> 11);
  assign _zz_mul_result_re_1 = ($signed(_zz_mul_result_re_2) - $signed(_zz_mul_result_re_3));
  assign _zz_mul_result_re_2 = ($signed(sub_result_re) * $signed(wn_re));
  assign _zz_mul_result_re_3 = ($signed(sub_result_im) * $signed(wn_im));
  assign _zz_mul_result_im = (_zz_mul_result_im_1 >>> 11);
  assign _zz_mul_result_im_1 = ($signed(_zz_mul_result_im_2) + $signed(_zz_mul_result_im_3));
  assign _zz_mul_result_im_2 = ($signed(sub_result_re) * $signed(wn_im));
  assign _zz_mul_result_im_3 = ($signed(sub_result_im) * $signed(wn_re));
  assign add_result_re = ($signed(in1_re) + $signed(in2_re));
  assign add_result_im = ($signed(in1_im) + $signed(in2_im));
  assign sub_result_re = ($signed(in1_re) - $signed(in2_re));
  assign sub_result_im = ($signed(in1_im) - $signed(in2_im));
  assign mul_result_re = _zz_mul_result_re[23:0];
  assign mul_result_im = _zz_mul_result_im[23:0];
  assign out1_re = add_result_re;
  assign out1_im = add_result_im;
  assign out2_re = mul_result_re;
  assign out2_im = mul_result_im;

endmodule

module ShiftRegisterNE (
  input      [23:0]   input_re,
  input      [23:0]   input_im,
  output     [23:0]   output_re,
  output     [23:0]   output_im,
  input               clk,
  input               reset
);
  reg        [23:0]   shift_reg_0_re;
  reg        [23:0]   shift_reg_0_im;
  reg        [23:0]   shift_reg_1_re;
  reg        [23:0]   shift_reg_1_im;
  reg        [23:0]   shift_reg_2_re;
  reg        [23:0]   shift_reg_2_im;
  reg        [23:0]   shift_reg_3_re;
  reg        [23:0]   shift_reg_3_im;
  reg        [23:0]   shift_reg_4_re;
  reg        [23:0]   shift_reg_4_im;
  reg        [23:0]   shift_reg_5_re;
  reg        [23:0]   shift_reg_5_im;
  reg        [23:0]   shift_reg_6_re;
  reg        [23:0]   shift_reg_6_im;
  reg        [23:0]   shift_reg_7_re;
  reg        [23:0]   shift_reg_7_im;
  reg        [23:0]   shift_reg_8_re;
  reg        [23:0]   shift_reg_8_im;
  reg        [23:0]   shift_reg_9_re;
  reg        [23:0]   shift_reg_9_im;
  reg        [23:0]   shift_reg_10_re;
  reg        [23:0]   shift_reg_10_im;
  reg        [23:0]   shift_reg_11_re;
  reg        [23:0]   shift_reg_11_im;
  reg        [23:0]   shift_reg_12_re;
  reg        [23:0]   shift_reg_12_im;
  reg        [23:0]   shift_reg_13_re;
  reg        [23:0]   shift_reg_13_im;
  reg        [23:0]   shift_reg_14_re;
  reg        [23:0]   shift_reg_14_im;
  reg        [23:0]   shift_reg_15_re;
  reg        [23:0]   shift_reg_15_im;
  reg        [23:0]   shift_reg_16_re;
  reg        [23:0]   shift_reg_16_im;
  reg        [23:0]   shift_reg_17_re;
  reg        [23:0]   shift_reg_17_im;
  reg        [23:0]   shift_reg_18_re;
  reg        [23:0]   shift_reg_18_im;
  reg        [23:0]   shift_reg_19_re;
  reg        [23:0]   shift_reg_19_im;
  reg        [23:0]   shift_reg_20_re;
  reg        [23:0]   shift_reg_20_im;
  reg        [23:0]   shift_reg_21_re;
  reg        [23:0]   shift_reg_21_im;
  reg        [23:0]   shift_reg_22_re;
  reg        [23:0]   shift_reg_22_im;
  reg        [23:0]   shift_reg_23_re;
  reg        [23:0]   shift_reg_23_im;
  reg        [23:0]   shift_reg_24_re;
  reg        [23:0]   shift_reg_24_im;
  reg        [23:0]   shift_reg_25_re;
  reg        [23:0]   shift_reg_25_im;
  reg        [23:0]   shift_reg_26_re;
  reg        [23:0]   shift_reg_26_im;
  reg        [23:0]   shift_reg_27_re;
  reg        [23:0]   shift_reg_27_im;
  reg        [23:0]   shift_reg_28_re;
  reg        [23:0]   shift_reg_28_im;
  reg        [23:0]   shift_reg_29_re;
  reg        [23:0]   shift_reg_29_im;
  reg        [23:0]   shift_reg_30_re;
  reg        [23:0]   shift_reg_30_im;
  reg        [23:0]   shift_reg_31_re;
  reg        [23:0]   shift_reg_31_im;
  reg        [23:0]   shift_reg_32_re;
  reg        [23:0]   shift_reg_32_im;
  reg        [23:0]   shift_reg_33_re;
  reg        [23:0]   shift_reg_33_im;
  reg        [23:0]   shift_reg_34_re;
  reg        [23:0]   shift_reg_34_im;
  reg        [23:0]   shift_reg_35_re;
  reg        [23:0]   shift_reg_35_im;
  reg        [23:0]   shift_reg_36_re;
  reg        [23:0]   shift_reg_36_im;
  reg        [23:0]   shift_reg_37_re;
  reg        [23:0]   shift_reg_37_im;
  reg        [23:0]   shift_reg_38_re;
  reg        [23:0]   shift_reg_38_im;
  reg        [23:0]   shift_reg_39_re;
  reg        [23:0]   shift_reg_39_im;
  reg        [23:0]   shift_reg_40_re;
  reg        [23:0]   shift_reg_40_im;
  reg        [23:0]   shift_reg_41_re;
  reg        [23:0]   shift_reg_41_im;
  reg        [23:0]   shift_reg_42_re;
  reg        [23:0]   shift_reg_42_im;
  reg        [23:0]   shift_reg_43_re;
  reg        [23:0]   shift_reg_43_im;
  reg        [23:0]   shift_reg_44_re;
  reg        [23:0]   shift_reg_44_im;
  reg        [23:0]   shift_reg_45_re;
  reg        [23:0]   shift_reg_45_im;
  reg        [23:0]   shift_reg_46_re;
  reg        [23:0]   shift_reg_46_im;
  reg        [23:0]   shift_reg_47_re;
  reg        [23:0]   shift_reg_47_im;
  reg        [23:0]   shift_reg_48_re;
  reg        [23:0]   shift_reg_48_im;
  reg        [23:0]   shift_reg_49_re;
  reg        [23:0]   shift_reg_49_im;
  reg        [23:0]   shift_reg_50_re;
  reg        [23:0]   shift_reg_50_im;
  reg        [23:0]   shift_reg_51_re;
  reg        [23:0]   shift_reg_51_im;
  reg        [23:0]   shift_reg_52_re;
  reg        [23:0]   shift_reg_52_im;
  reg        [23:0]   shift_reg_53_re;
  reg        [23:0]   shift_reg_53_im;
  reg        [23:0]   shift_reg_54_re;
  reg        [23:0]   shift_reg_54_im;
  reg        [23:0]   shift_reg_55_re;
  reg        [23:0]   shift_reg_55_im;
  reg        [23:0]   shift_reg_56_re;
  reg        [23:0]   shift_reg_56_im;
  reg        [23:0]   shift_reg_57_re;
  reg        [23:0]   shift_reg_57_im;
  reg        [23:0]   shift_reg_58_re;
  reg        [23:0]   shift_reg_58_im;
  reg        [23:0]   shift_reg_59_re;
  reg        [23:0]   shift_reg_59_im;
  reg        [23:0]   shift_reg_60_re;
  reg        [23:0]   shift_reg_60_im;
  reg        [23:0]   shift_reg_61_re;
  reg        [23:0]   shift_reg_61_im;
  reg        [23:0]   shift_reg_62_re;
  reg        [23:0]   shift_reg_62_im;
  reg        [23:0]   shift_reg_63_re;
  reg        [23:0]   shift_reg_63_im;
  reg        [23:0]   shift_reg_64_re;
  reg        [23:0]   shift_reg_64_im;
  reg        [23:0]   shift_reg_65_re;
  reg        [23:0]   shift_reg_65_im;
  reg        [23:0]   shift_reg_66_re;
  reg        [23:0]   shift_reg_66_im;
  reg        [23:0]   shift_reg_67_re;
  reg        [23:0]   shift_reg_67_im;
  reg        [23:0]   shift_reg_68_re;
  reg        [23:0]   shift_reg_68_im;
  reg        [23:0]   shift_reg_69_re;
  reg        [23:0]   shift_reg_69_im;
  reg        [23:0]   shift_reg_70_re;
  reg        [23:0]   shift_reg_70_im;
  reg        [23:0]   shift_reg_71_re;
  reg        [23:0]   shift_reg_71_im;
  reg        [23:0]   shift_reg_72_re;
  reg        [23:0]   shift_reg_72_im;
  reg        [23:0]   shift_reg_73_re;
  reg        [23:0]   shift_reg_73_im;
  reg        [23:0]   shift_reg_74_re;
  reg        [23:0]   shift_reg_74_im;
  reg        [23:0]   shift_reg_75_re;
  reg        [23:0]   shift_reg_75_im;
  reg        [23:0]   shift_reg_76_re;
  reg        [23:0]   shift_reg_76_im;
  reg        [23:0]   shift_reg_77_re;
  reg        [23:0]   shift_reg_77_im;
  reg        [23:0]   shift_reg_78_re;
  reg        [23:0]   shift_reg_78_im;
  reg        [23:0]   shift_reg_79_re;
  reg        [23:0]   shift_reg_79_im;
  reg        [23:0]   shift_reg_80_re;
  reg        [23:0]   shift_reg_80_im;
  reg        [23:0]   shift_reg_81_re;
  reg        [23:0]   shift_reg_81_im;
  reg        [23:0]   shift_reg_82_re;
  reg        [23:0]   shift_reg_82_im;
  reg        [23:0]   shift_reg_83_re;
  reg        [23:0]   shift_reg_83_im;
  reg        [23:0]   shift_reg_84_re;
  reg        [23:0]   shift_reg_84_im;
  reg        [23:0]   shift_reg_85_re;
  reg        [23:0]   shift_reg_85_im;
  reg        [23:0]   shift_reg_86_re;
  reg        [23:0]   shift_reg_86_im;
  reg        [23:0]   shift_reg_87_re;
  reg        [23:0]   shift_reg_87_im;
  reg        [23:0]   shift_reg_88_re;
  reg        [23:0]   shift_reg_88_im;
  reg        [23:0]   shift_reg_89_re;
  reg        [23:0]   shift_reg_89_im;
  reg        [23:0]   shift_reg_90_re;
  reg        [23:0]   shift_reg_90_im;
  reg        [23:0]   shift_reg_91_re;
  reg        [23:0]   shift_reg_91_im;
  reg        [23:0]   shift_reg_92_re;
  reg        [23:0]   shift_reg_92_im;
  reg        [23:0]   shift_reg_93_re;
  reg        [23:0]   shift_reg_93_im;
  reg        [23:0]   shift_reg_94_re;
  reg        [23:0]   shift_reg_94_im;
  reg        [23:0]   shift_reg_95_re;
  reg        [23:0]   shift_reg_95_im;
  reg        [23:0]   shift_reg_96_re;
  reg        [23:0]   shift_reg_96_im;
  reg        [23:0]   shift_reg_97_re;
  reg        [23:0]   shift_reg_97_im;
  reg        [23:0]   shift_reg_98_re;
  reg        [23:0]   shift_reg_98_im;
  reg        [23:0]   shift_reg_99_re;
  reg        [23:0]   shift_reg_99_im;
  reg        [23:0]   shift_reg_100_re;
  reg        [23:0]   shift_reg_100_im;
  reg        [23:0]   shift_reg_101_re;
  reg        [23:0]   shift_reg_101_im;
  reg        [23:0]   shift_reg_102_re;
  reg        [23:0]   shift_reg_102_im;
  reg        [23:0]   shift_reg_103_re;
  reg        [23:0]   shift_reg_103_im;
  reg        [23:0]   shift_reg_104_re;
  reg        [23:0]   shift_reg_104_im;
  reg        [23:0]   shift_reg_105_re;
  reg        [23:0]   shift_reg_105_im;
  reg        [23:0]   shift_reg_106_re;
  reg        [23:0]   shift_reg_106_im;
  reg        [23:0]   shift_reg_107_re;
  reg        [23:0]   shift_reg_107_im;
  reg        [23:0]   shift_reg_108_re;
  reg        [23:0]   shift_reg_108_im;
  reg        [23:0]   shift_reg_109_re;
  reg        [23:0]   shift_reg_109_im;
  reg        [23:0]   shift_reg_110_re;
  reg        [23:0]   shift_reg_110_im;
  reg        [23:0]   shift_reg_111_re;
  reg        [23:0]   shift_reg_111_im;
  reg        [23:0]   shift_reg_112_re;
  reg        [23:0]   shift_reg_112_im;
  reg        [23:0]   shift_reg_113_re;
  reg        [23:0]   shift_reg_113_im;
  reg        [23:0]   shift_reg_114_re;
  reg        [23:0]   shift_reg_114_im;
  reg        [23:0]   shift_reg_115_re;
  reg        [23:0]   shift_reg_115_im;
  reg        [23:0]   shift_reg_116_re;
  reg        [23:0]   shift_reg_116_im;
  reg        [23:0]   shift_reg_117_re;
  reg        [23:0]   shift_reg_117_im;
  reg        [23:0]   shift_reg_118_re;
  reg        [23:0]   shift_reg_118_im;
  reg        [23:0]   shift_reg_119_re;
  reg        [23:0]   shift_reg_119_im;
  reg        [23:0]   shift_reg_120_re;
  reg        [23:0]   shift_reg_120_im;
  reg        [23:0]   shift_reg_121_re;
  reg        [23:0]   shift_reg_121_im;
  reg        [23:0]   shift_reg_122_re;
  reg        [23:0]   shift_reg_122_im;
  reg        [23:0]   shift_reg_123_re;
  reg        [23:0]   shift_reg_123_im;
  reg        [23:0]   shift_reg_124_re;
  reg        [23:0]   shift_reg_124_im;
  reg        [23:0]   shift_reg_125_re;
  reg        [23:0]   shift_reg_125_im;
  reg        [23:0]   shift_reg_126_re;
  reg        [23:0]   shift_reg_126_im;
  reg        [23:0]   shift_reg_127_re;
  reg        [23:0]   shift_reg_127_im;
  reg        [23:0]   shift_reg_128_re;
  reg        [23:0]   shift_reg_128_im;
  reg        [23:0]   shift_reg_129_re;
  reg        [23:0]   shift_reg_129_im;
  reg        [23:0]   shift_reg_130_re;
  reg        [23:0]   shift_reg_130_im;
  reg        [23:0]   shift_reg_131_re;
  reg        [23:0]   shift_reg_131_im;
  reg        [23:0]   shift_reg_132_re;
  reg        [23:0]   shift_reg_132_im;
  reg        [23:0]   shift_reg_133_re;
  reg        [23:0]   shift_reg_133_im;
  reg        [23:0]   shift_reg_134_re;
  reg        [23:0]   shift_reg_134_im;
  reg        [23:0]   shift_reg_135_re;
  reg        [23:0]   shift_reg_135_im;
  reg        [23:0]   shift_reg_136_re;
  reg        [23:0]   shift_reg_136_im;
  reg        [23:0]   shift_reg_137_re;
  reg        [23:0]   shift_reg_137_im;
  reg        [23:0]   shift_reg_138_re;
  reg        [23:0]   shift_reg_138_im;
  reg        [23:0]   shift_reg_139_re;
  reg        [23:0]   shift_reg_139_im;
  reg        [23:0]   shift_reg_140_re;
  reg        [23:0]   shift_reg_140_im;
  reg        [23:0]   shift_reg_141_re;
  reg        [23:0]   shift_reg_141_im;
  reg        [23:0]   shift_reg_142_re;
  reg        [23:0]   shift_reg_142_im;
  reg        [23:0]   shift_reg_143_re;
  reg        [23:0]   shift_reg_143_im;
  reg        [23:0]   shift_reg_144_re;
  reg        [23:0]   shift_reg_144_im;
  reg        [23:0]   shift_reg_145_re;
  reg        [23:0]   shift_reg_145_im;
  reg        [23:0]   shift_reg_146_re;
  reg        [23:0]   shift_reg_146_im;
  reg        [23:0]   shift_reg_147_re;
  reg        [23:0]   shift_reg_147_im;
  reg        [23:0]   shift_reg_148_re;
  reg        [23:0]   shift_reg_148_im;
  reg        [23:0]   shift_reg_149_re;
  reg        [23:0]   shift_reg_149_im;
  reg        [23:0]   shift_reg_150_re;
  reg        [23:0]   shift_reg_150_im;
  reg        [23:0]   shift_reg_151_re;
  reg        [23:0]   shift_reg_151_im;
  reg        [23:0]   shift_reg_152_re;
  reg        [23:0]   shift_reg_152_im;
  reg        [23:0]   shift_reg_153_re;
  reg        [23:0]   shift_reg_153_im;
  reg        [23:0]   shift_reg_154_re;
  reg        [23:0]   shift_reg_154_im;
  reg        [23:0]   shift_reg_155_re;
  reg        [23:0]   shift_reg_155_im;
  reg        [23:0]   shift_reg_156_re;
  reg        [23:0]   shift_reg_156_im;
  reg        [23:0]   shift_reg_157_re;
  reg        [23:0]   shift_reg_157_im;
  reg        [23:0]   shift_reg_158_re;
  reg        [23:0]   shift_reg_158_im;
  reg        [23:0]   shift_reg_159_re;
  reg        [23:0]   shift_reg_159_im;
  reg        [23:0]   shift_reg_160_re;
  reg        [23:0]   shift_reg_160_im;
  reg        [23:0]   shift_reg_161_re;
  reg        [23:0]   shift_reg_161_im;
  reg        [23:0]   shift_reg_162_re;
  reg        [23:0]   shift_reg_162_im;
  reg        [23:0]   shift_reg_163_re;
  reg        [23:0]   shift_reg_163_im;
  reg        [23:0]   shift_reg_164_re;
  reg        [23:0]   shift_reg_164_im;
  reg        [23:0]   shift_reg_165_re;
  reg        [23:0]   shift_reg_165_im;
  reg        [23:0]   shift_reg_166_re;
  reg        [23:0]   shift_reg_166_im;
  reg        [23:0]   shift_reg_167_re;
  reg        [23:0]   shift_reg_167_im;
  reg        [23:0]   shift_reg_168_re;
  reg        [23:0]   shift_reg_168_im;
  reg        [23:0]   shift_reg_169_re;
  reg        [23:0]   shift_reg_169_im;
  reg        [23:0]   shift_reg_170_re;
  reg        [23:0]   shift_reg_170_im;
  reg        [23:0]   shift_reg_171_re;
  reg        [23:0]   shift_reg_171_im;
  reg        [23:0]   shift_reg_172_re;
  reg        [23:0]   shift_reg_172_im;
  reg        [23:0]   shift_reg_173_re;
  reg        [23:0]   shift_reg_173_im;
  reg        [23:0]   shift_reg_174_re;
  reg        [23:0]   shift_reg_174_im;
  reg        [23:0]   shift_reg_175_re;
  reg        [23:0]   shift_reg_175_im;
  reg        [23:0]   shift_reg_176_re;
  reg        [23:0]   shift_reg_176_im;
  reg        [23:0]   shift_reg_177_re;
  reg        [23:0]   shift_reg_177_im;
  reg        [23:0]   shift_reg_178_re;
  reg        [23:0]   shift_reg_178_im;
  reg        [23:0]   shift_reg_179_re;
  reg        [23:0]   shift_reg_179_im;
  reg        [23:0]   shift_reg_180_re;
  reg        [23:0]   shift_reg_180_im;
  reg        [23:0]   shift_reg_181_re;
  reg        [23:0]   shift_reg_181_im;
  reg        [23:0]   shift_reg_182_re;
  reg        [23:0]   shift_reg_182_im;
  reg        [23:0]   shift_reg_183_re;
  reg        [23:0]   shift_reg_183_im;
  reg        [23:0]   shift_reg_184_re;
  reg        [23:0]   shift_reg_184_im;
  reg        [23:0]   shift_reg_185_re;
  reg        [23:0]   shift_reg_185_im;
  reg        [23:0]   shift_reg_186_re;
  reg        [23:0]   shift_reg_186_im;
  reg        [23:0]   shift_reg_187_re;
  reg        [23:0]   shift_reg_187_im;
  reg        [23:0]   shift_reg_188_re;
  reg        [23:0]   shift_reg_188_im;
  reg        [23:0]   shift_reg_189_re;
  reg        [23:0]   shift_reg_189_im;
  reg        [23:0]   shift_reg_190_re;
  reg        [23:0]   shift_reg_190_im;
  reg        [23:0]   shift_reg_191_re;
  reg        [23:0]   shift_reg_191_im;
  reg        [23:0]   shift_reg_192_re;
  reg        [23:0]   shift_reg_192_im;
  reg        [23:0]   shift_reg_193_re;
  reg        [23:0]   shift_reg_193_im;
  reg        [23:0]   shift_reg_194_re;
  reg        [23:0]   shift_reg_194_im;
  reg        [23:0]   shift_reg_195_re;
  reg        [23:0]   shift_reg_195_im;
  reg        [23:0]   shift_reg_196_re;
  reg        [23:0]   shift_reg_196_im;
  reg        [23:0]   shift_reg_197_re;
  reg        [23:0]   shift_reg_197_im;
  reg        [23:0]   shift_reg_198_re;
  reg        [23:0]   shift_reg_198_im;
  reg        [23:0]   shift_reg_199_re;
  reg        [23:0]   shift_reg_199_im;
  reg        [23:0]   shift_reg_200_re;
  reg        [23:0]   shift_reg_200_im;
  reg        [23:0]   shift_reg_201_re;
  reg        [23:0]   shift_reg_201_im;
  reg        [23:0]   shift_reg_202_re;
  reg        [23:0]   shift_reg_202_im;
  reg        [23:0]   shift_reg_203_re;
  reg        [23:0]   shift_reg_203_im;
  reg        [23:0]   shift_reg_204_re;
  reg        [23:0]   shift_reg_204_im;
  reg        [23:0]   shift_reg_205_re;
  reg        [23:0]   shift_reg_205_im;
  reg        [23:0]   shift_reg_206_re;
  reg        [23:0]   shift_reg_206_im;
  reg        [23:0]   shift_reg_207_re;
  reg        [23:0]   shift_reg_207_im;
  reg        [23:0]   shift_reg_208_re;
  reg        [23:0]   shift_reg_208_im;
  reg        [23:0]   shift_reg_209_re;
  reg        [23:0]   shift_reg_209_im;
  reg        [23:0]   shift_reg_210_re;
  reg        [23:0]   shift_reg_210_im;
  reg        [23:0]   shift_reg_211_re;
  reg        [23:0]   shift_reg_211_im;
  reg        [23:0]   shift_reg_212_re;
  reg        [23:0]   shift_reg_212_im;
  reg        [23:0]   shift_reg_213_re;
  reg        [23:0]   shift_reg_213_im;
  reg        [23:0]   shift_reg_214_re;
  reg        [23:0]   shift_reg_214_im;
  reg        [23:0]   shift_reg_215_re;
  reg        [23:0]   shift_reg_215_im;
  reg        [23:0]   shift_reg_216_re;
  reg        [23:0]   shift_reg_216_im;
  reg        [23:0]   shift_reg_217_re;
  reg        [23:0]   shift_reg_217_im;
  reg        [23:0]   shift_reg_218_re;
  reg        [23:0]   shift_reg_218_im;
  reg        [23:0]   shift_reg_219_re;
  reg        [23:0]   shift_reg_219_im;
  reg        [23:0]   shift_reg_220_re;
  reg        [23:0]   shift_reg_220_im;
  reg        [23:0]   shift_reg_221_re;
  reg        [23:0]   shift_reg_221_im;
  reg        [23:0]   shift_reg_222_re;
  reg        [23:0]   shift_reg_222_im;
  reg        [23:0]   shift_reg_223_re;
  reg        [23:0]   shift_reg_223_im;
  reg        [23:0]   shift_reg_224_re;
  reg        [23:0]   shift_reg_224_im;
  reg        [23:0]   shift_reg_225_re;
  reg        [23:0]   shift_reg_225_im;
  reg        [23:0]   shift_reg_226_re;
  reg        [23:0]   shift_reg_226_im;
  reg        [23:0]   shift_reg_227_re;
  reg        [23:0]   shift_reg_227_im;
  reg        [23:0]   shift_reg_228_re;
  reg        [23:0]   shift_reg_228_im;
  reg        [23:0]   shift_reg_229_re;
  reg        [23:0]   shift_reg_229_im;
  reg        [23:0]   shift_reg_230_re;
  reg        [23:0]   shift_reg_230_im;
  reg        [23:0]   shift_reg_231_re;
  reg        [23:0]   shift_reg_231_im;
  reg        [23:0]   shift_reg_232_re;
  reg        [23:0]   shift_reg_232_im;
  reg        [23:0]   shift_reg_233_re;
  reg        [23:0]   shift_reg_233_im;
  reg        [23:0]   shift_reg_234_re;
  reg        [23:0]   shift_reg_234_im;
  reg        [23:0]   shift_reg_235_re;
  reg        [23:0]   shift_reg_235_im;
  reg        [23:0]   shift_reg_236_re;
  reg        [23:0]   shift_reg_236_im;
  reg        [23:0]   shift_reg_237_re;
  reg        [23:0]   shift_reg_237_im;
  reg        [23:0]   shift_reg_238_re;
  reg        [23:0]   shift_reg_238_im;
  reg        [23:0]   shift_reg_239_re;
  reg        [23:0]   shift_reg_239_im;
  reg        [23:0]   shift_reg_240_re;
  reg        [23:0]   shift_reg_240_im;
  reg        [23:0]   shift_reg_241_re;
  reg        [23:0]   shift_reg_241_im;
  reg        [23:0]   shift_reg_242_re;
  reg        [23:0]   shift_reg_242_im;
  reg        [23:0]   shift_reg_243_re;
  reg        [23:0]   shift_reg_243_im;
  reg        [23:0]   shift_reg_244_re;
  reg        [23:0]   shift_reg_244_im;
  reg        [23:0]   shift_reg_245_re;
  reg        [23:0]   shift_reg_245_im;
  reg        [23:0]   shift_reg_246_re;
  reg        [23:0]   shift_reg_246_im;
  reg        [23:0]   shift_reg_247_re;
  reg        [23:0]   shift_reg_247_im;
  reg        [23:0]   shift_reg_248_re;
  reg        [23:0]   shift_reg_248_im;
  reg        [23:0]   shift_reg_249_re;
  reg        [23:0]   shift_reg_249_im;
  reg        [23:0]   shift_reg_250_re;
  reg        [23:0]   shift_reg_250_im;
  reg        [23:0]   shift_reg_251_re;
  reg        [23:0]   shift_reg_251_im;
  reg        [23:0]   shift_reg_252_re;
  reg        [23:0]   shift_reg_252_im;
  reg        [23:0]   shift_reg_253_re;
  reg        [23:0]   shift_reg_253_im;
  reg        [23:0]   shift_reg_254_re;
  reg        [23:0]   shift_reg_254_im;
  reg        [23:0]   shift_reg_255_re;
  reg        [23:0]   shift_reg_255_im;
  reg        [23:0]   shift_reg_256_re;
  reg        [23:0]   shift_reg_256_im;
  reg        [23:0]   shift_reg_257_re;
  reg        [23:0]   shift_reg_257_im;
  reg        [23:0]   shift_reg_258_re;
  reg        [23:0]   shift_reg_258_im;
  reg        [23:0]   shift_reg_259_re;
  reg        [23:0]   shift_reg_259_im;
  reg        [23:0]   shift_reg_260_re;
  reg        [23:0]   shift_reg_260_im;
  reg        [23:0]   shift_reg_261_re;
  reg        [23:0]   shift_reg_261_im;
  reg        [23:0]   shift_reg_262_re;
  reg        [23:0]   shift_reg_262_im;
  reg        [23:0]   shift_reg_263_re;
  reg        [23:0]   shift_reg_263_im;
  reg        [23:0]   shift_reg_264_re;
  reg        [23:0]   shift_reg_264_im;
  reg        [23:0]   shift_reg_265_re;
  reg        [23:0]   shift_reg_265_im;
  reg        [23:0]   shift_reg_266_re;
  reg        [23:0]   shift_reg_266_im;
  reg        [23:0]   shift_reg_267_re;
  reg        [23:0]   shift_reg_267_im;
  reg        [23:0]   shift_reg_268_re;
  reg        [23:0]   shift_reg_268_im;
  reg        [23:0]   shift_reg_269_re;
  reg        [23:0]   shift_reg_269_im;
  reg        [23:0]   shift_reg_270_re;
  reg        [23:0]   shift_reg_270_im;
  reg        [23:0]   shift_reg_271_re;
  reg        [23:0]   shift_reg_271_im;
  reg        [23:0]   shift_reg_272_re;
  reg        [23:0]   shift_reg_272_im;
  reg        [23:0]   shift_reg_273_re;
  reg        [23:0]   shift_reg_273_im;
  reg        [23:0]   shift_reg_274_re;
  reg        [23:0]   shift_reg_274_im;
  reg        [23:0]   shift_reg_275_re;
  reg        [23:0]   shift_reg_275_im;
  reg        [23:0]   shift_reg_276_re;
  reg        [23:0]   shift_reg_276_im;
  reg        [23:0]   shift_reg_277_re;
  reg        [23:0]   shift_reg_277_im;
  reg        [23:0]   shift_reg_278_re;
  reg        [23:0]   shift_reg_278_im;
  reg        [23:0]   shift_reg_279_re;
  reg        [23:0]   shift_reg_279_im;
  reg        [23:0]   shift_reg_280_re;
  reg        [23:0]   shift_reg_280_im;
  reg        [23:0]   shift_reg_281_re;
  reg        [23:0]   shift_reg_281_im;
  reg        [23:0]   shift_reg_282_re;
  reg        [23:0]   shift_reg_282_im;
  reg        [23:0]   shift_reg_283_re;
  reg        [23:0]   shift_reg_283_im;
  reg        [23:0]   shift_reg_284_re;
  reg        [23:0]   shift_reg_284_im;
  reg        [23:0]   shift_reg_285_re;
  reg        [23:0]   shift_reg_285_im;
  reg        [23:0]   shift_reg_286_re;
  reg        [23:0]   shift_reg_286_im;
  reg        [23:0]   shift_reg_287_re;
  reg        [23:0]   shift_reg_287_im;
  reg        [23:0]   shift_reg_288_re;
  reg        [23:0]   shift_reg_288_im;
  reg        [23:0]   shift_reg_289_re;
  reg        [23:0]   shift_reg_289_im;
  reg        [23:0]   shift_reg_290_re;
  reg        [23:0]   shift_reg_290_im;
  reg        [23:0]   shift_reg_291_re;
  reg        [23:0]   shift_reg_291_im;
  reg        [23:0]   shift_reg_292_re;
  reg        [23:0]   shift_reg_292_im;
  reg        [23:0]   shift_reg_293_re;
  reg        [23:0]   shift_reg_293_im;
  reg        [23:0]   shift_reg_294_re;
  reg        [23:0]   shift_reg_294_im;
  reg        [23:0]   shift_reg_295_re;
  reg        [23:0]   shift_reg_295_im;
  reg        [23:0]   shift_reg_296_re;
  reg        [23:0]   shift_reg_296_im;
  reg        [23:0]   shift_reg_297_re;
  reg        [23:0]   shift_reg_297_im;
  reg        [23:0]   shift_reg_298_re;
  reg        [23:0]   shift_reg_298_im;
  reg        [23:0]   shift_reg_299_re;
  reg        [23:0]   shift_reg_299_im;
  reg        [23:0]   shift_reg_300_re;
  reg        [23:0]   shift_reg_300_im;
  reg        [23:0]   shift_reg_301_re;
  reg        [23:0]   shift_reg_301_im;
  reg        [23:0]   shift_reg_302_re;
  reg        [23:0]   shift_reg_302_im;
  reg        [23:0]   shift_reg_303_re;
  reg        [23:0]   shift_reg_303_im;
  reg        [23:0]   shift_reg_304_re;
  reg        [23:0]   shift_reg_304_im;
  reg        [23:0]   shift_reg_305_re;
  reg        [23:0]   shift_reg_305_im;
  reg        [23:0]   shift_reg_306_re;
  reg        [23:0]   shift_reg_306_im;
  reg        [23:0]   shift_reg_307_re;
  reg        [23:0]   shift_reg_307_im;
  reg        [23:0]   shift_reg_308_re;
  reg        [23:0]   shift_reg_308_im;
  reg        [23:0]   shift_reg_309_re;
  reg        [23:0]   shift_reg_309_im;
  reg        [23:0]   shift_reg_310_re;
  reg        [23:0]   shift_reg_310_im;
  reg        [23:0]   shift_reg_311_re;
  reg        [23:0]   shift_reg_311_im;
  reg        [23:0]   shift_reg_312_re;
  reg        [23:0]   shift_reg_312_im;
  reg        [23:0]   shift_reg_313_re;
  reg        [23:0]   shift_reg_313_im;
  reg        [23:0]   shift_reg_314_re;
  reg        [23:0]   shift_reg_314_im;
  reg        [23:0]   shift_reg_315_re;
  reg        [23:0]   shift_reg_315_im;
  reg        [23:0]   shift_reg_316_re;
  reg        [23:0]   shift_reg_316_im;
  reg        [23:0]   shift_reg_317_re;
  reg        [23:0]   shift_reg_317_im;
  reg        [23:0]   shift_reg_318_re;
  reg        [23:0]   shift_reg_318_im;
  reg        [23:0]   shift_reg_319_re;
  reg        [23:0]   shift_reg_319_im;
  reg        [23:0]   shift_reg_320_re;
  reg        [23:0]   shift_reg_320_im;
  reg        [23:0]   shift_reg_321_re;
  reg        [23:0]   shift_reg_321_im;
  reg        [23:0]   shift_reg_322_re;
  reg        [23:0]   shift_reg_322_im;
  reg        [23:0]   shift_reg_323_re;
  reg        [23:0]   shift_reg_323_im;
  reg        [23:0]   shift_reg_324_re;
  reg        [23:0]   shift_reg_324_im;
  reg        [23:0]   shift_reg_325_re;
  reg        [23:0]   shift_reg_325_im;
  reg        [23:0]   shift_reg_326_re;
  reg        [23:0]   shift_reg_326_im;
  reg        [23:0]   shift_reg_327_re;
  reg        [23:0]   shift_reg_327_im;
  reg        [23:0]   shift_reg_328_re;
  reg        [23:0]   shift_reg_328_im;
  reg        [23:0]   shift_reg_329_re;
  reg        [23:0]   shift_reg_329_im;
  reg        [23:0]   shift_reg_330_re;
  reg        [23:0]   shift_reg_330_im;
  reg        [23:0]   shift_reg_331_re;
  reg        [23:0]   shift_reg_331_im;
  reg        [23:0]   shift_reg_332_re;
  reg        [23:0]   shift_reg_332_im;
  reg        [23:0]   shift_reg_333_re;
  reg        [23:0]   shift_reg_333_im;
  reg        [23:0]   shift_reg_334_re;
  reg        [23:0]   shift_reg_334_im;
  reg        [23:0]   shift_reg_335_re;
  reg        [23:0]   shift_reg_335_im;
  reg        [23:0]   shift_reg_336_re;
  reg        [23:0]   shift_reg_336_im;
  reg        [23:0]   shift_reg_337_re;
  reg        [23:0]   shift_reg_337_im;
  reg        [23:0]   shift_reg_338_re;
  reg        [23:0]   shift_reg_338_im;
  reg        [23:0]   shift_reg_339_re;
  reg        [23:0]   shift_reg_339_im;
  reg        [23:0]   shift_reg_340_re;
  reg        [23:0]   shift_reg_340_im;
  reg        [23:0]   shift_reg_341_re;
  reg        [23:0]   shift_reg_341_im;
  reg        [23:0]   shift_reg_342_re;
  reg        [23:0]   shift_reg_342_im;
  reg        [23:0]   shift_reg_343_re;
  reg        [23:0]   shift_reg_343_im;
  reg        [23:0]   shift_reg_344_re;
  reg        [23:0]   shift_reg_344_im;
  reg        [23:0]   shift_reg_345_re;
  reg        [23:0]   shift_reg_345_im;
  reg        [23:0]   shift_reg_346_re;
  reg        [23:0]   shift_reg_346_im;
  reg        [23:0]   shift_reg_347_re;
  reg        [23:0]   shift_reg_347_im;
  reg        [23:0]   shift_reg_348_re;
  reg        [23:0]   shift_reg_348_im;
  reg        [23:0]   shift_reg_349_re;
  reg        [23:0]   shift_reg_349_im;
  reg        [23:0]   shift_reg_350_re;
  reg        [23:0]   shift_reg_350_im;
  reg        [23:0]   shift_reg_351_re;
  reg        [23:0]   shift_reg_351_im;
  reg        [23:0]   shift_reg_352_re;
  reg        [23:0]   shift_reg_352_im;
  reg        [23:0]   shift_reg_353_re;
  reg        [23:0]   shift_reg_353_im;
  reg        [23:0]   shift_reg_354_re;
  reg        [23:0]   shift_reg_354_im;
  reg        [23:0]   shift_reg_355_re;
  reg        [23:0]   shift_reg_355_im;
  reg        [23:0]   shift_reg_356_re;
  reg        [23:0]   shift_reg_356_im;
  reg        [23:0]   shift_reg_357_re;
  reg        [23:0]   shift_reg_357_im;
  reg        [23:0]   shift_reg_358_re;
  reg        [23:0]   shift_reg_358_im;
  reg        [23:0]   shift_reg_359_re;
  reg        [23:0]   shift_reg_359_im;
  reg        [23:0]   shift_reg_360_re;
  reg        [23:0]   shift_reg_360_im;
  reg        [23:0]   shift_reg_361_re;
  reg        [23:0]   shift_reg_361_im;
  reg        [23:0]   shift_reg_362_re;
  reg        [23:0]   shift_reg_362_im;
  reg        [23:0]   shift_reg_363_re;
  reg        [23:0]   shift_reg_363_im;
  reg        [23:0]   shift_reg_364_re;
  reg        [23:0]   shift_reg_364_im;
  reg        [23:0]   shift_reg_365_re;
  reg        [23:0]   shift_reg_365_im;
  reg        [23:0]   shift_reg_366_re;
  reg        [23:0]   shift_reg_366_im;
  reg        [23:0]   shift_reg_367_re;
  reg        [23:0]   shift_reg_367_im;
  reg        [23:0]   shift_reg_368_re;
  reg        [23:0]   shift_reg_368_im;
  reg        [23:0]   shift_reg_369_re;
  reg        [23:0]   shift_reg_369_im;
  reg        [23:0]   shift_reg_370_re;
  reg        [23:0]   shift_reg_370_im;
  reg        [23:0]   shift_reg_371_re;
  reg        [23:0]   shift_reg_371_im;
  reg        [23:0]   shift_reg_372_re;
  reg        [23:0]   shift_reg_372_im;
  reg        [23:0]   shift_reg_373_re;
  reg        [23:0]   shift_reg_373_im;
  reg        [23:0]   shift_reg_374_re;
  reg        [23:0]   shift_reg_374_im;
  reg        [23:0]   shift_reg_375_re;
  reg        [23:0]   shift_reg_375_im;
  reg        [23:0]   shift_reg_376_re;
  reg        [23:0]   shift_reg_376_im;
  reg        [23:0]   shift_reg_377_re;
  reg        [23:0]   shift_reg_377_im;
  reg        [23:0]   shift_reg_378_re;
  reg        [23:0]   shift_reg_378_im;
  reg        [23:0]   shift_reg_379_re;
  reg        [23:0]   shift_reg_379_im;
  reg        [23:0]   shift_reg_380_re;
  reg        [23:0]   shift_reg_380_im;
  reg        [23:0]   shift_reg_381_re;
  reg        [23:0]   shift_reg_381_im;
  reg        [23:0]   shift_reg_382_re;
  reg        [23:0]   shift_reg_382_im;
  reg        [23:0]   shift_reg_383_re;
  reg        [23:0]   shift_reg_383_im;
  reg        [23:0]   shift_reg_384_re;
  reg        [23:0]   shift_reg_384_im;
  reg        [23:0]   shift_reg_385_re;
  reg        [23:0]   shift_reg_385_im;
  reg        [23:0]   shift_reg_386_re;
  reg        [23:0]   shift_reg_386_im;
  reg        [23:0]   shift_reg_387_re;
  reg        [23:0]   shift_reg_387_im;
  reg        [23:0]   shift_reg_388_re;
  reg        [23:0]   shift_reg_388_im;
  reg        [23:0]   shift_reg_389_re;
  reg        [23:0]   shift_reg_389_im;
  reg        [23:0]   shift_reg_390_re;
  reg        [23:0]   shift_reg_390_im;
  reg        [23:0]   shift_reg_391_re;
  reg        [23:0]   shift_reg_391_im;
  reg        [23:0]   shift_reg_392_re;
  reg        [23:0]   shift_reg_392_im;
  reg        [23:0]   shift_reg_393_re;
  reg        [23:0]   shift_reg_393_im;
  reg        [23:0]   shift_reg_394_re;
  reg        [23:0]   shift_reg_394_im;
  reg        [23:0]   shift_reg_395_re;
  reg        [23:0]   shift_reg_395_im;
  reg        [23:0]   shift_reg_396_re;
  reg        [23:0]   shift_reg_396_im;
  reg        [23:0]   shift_reg_397_re;
  reg        [23:0]   shift_reg_397_im;
  reg        [23:0]   shift_reg_398_re;
  reg        [23:0]   shift_reg_398_im;
  reg        [23:0]   shift_reg_399_re;
  reg        [23:0]   shift_reg_399_im;
  reg        [23:0]   shift_reg_400_re;
  reg        [23:0]   shift_reg_400_im;
  reg        [23:0]   shift_reg_401_re;
  reg        [23:0]   shift_reg_401_im;
  reg        [23:0]   shift_reg_402_re;
  reg        [23:0]   shift_reg_402_im;
  reg        [23:0]   shift_reg_403_re;
  reg        [23:0]   shift_reg_403_im;
  reg        [23:0]   shift_reg_404_re;
  reg        [23:0]   shift_reg_404_im;
  reg        [23:0]   shift_reg_405_re;
  reg        [23:0]   shift_reg_405_im;
  reg        [23:0]   shift_reg_406_re;
  reg        [23:0]   shift_reg_406_im;
  reg        [23:0]   shift_reg_407_re;
  reg        [23:0]   shift_reg_407_im;
  reg        [23:0]   shift_reg_408_re;
  reg        [23:0]   shift_reg_408_im;
  reg        [23:0]   shift_reg_409_re;
  reg        [23:0]   shift_reg_409_im;
  reg        [23:0]   shift_reg_410_re;
  reg        [23:0]   shift_reg_410_im;
  reg        [23:0]   shift_reg_411_re;
  reg        [23:0]   shift_reg_411_im;
  reg        [23:0]   shift_reg_412_re;
  reg        [23:0]   shift_reg_412_im;
  reg        [23:0]   shift_reg_413_re;
  reg        [23:0]   shift_reg_413_im;
  reg        [23:0]   shift_reg_414_re;
  reg        [23:0]   shift_reg_414_im;
  reg        [23:0]   shift_reg_415_re;
  reg        [23:0]   shift_reg_415_im;
  reg        [23:0]   shift_reg_416_re;
  reg        [23:0]   shift_reg_416_im;
  reg        [23:0]   shift_reg_417_re;
  reg        [23:0]   shift_reg_417_im;
  reg        [23:0]   shift_reg_418_re;
  reg        [23:0]   shift_reg_418_im;
  reg        [23:0]   shift_reg_419_re;
  reg        [23:0]   shift_reg_419_im;
  reg        [23:0]   shift_reg_420_re;
  reg        [23:0]   shift_reg_420_im;
  reg        [23:0]   shift_reg_421_re;
  reg        [23:0]   shift_reg_421_im;
  reg        [23:0]   shift_reg_422_re;
  reg        [23:0]   shift_reg_422_im;
  reg        [23:0]   shift_reg_423_re;
  reg        [23:0]   shift_reg_423_im;
  reg        [23:0]   shift_reg_424_re;
  reg        [23:0]   shift_reg_424_im;
  reg        [23:0]   shift_reg_425_re;
  reg        [23:0]   shift_reg_425_im;
  reg        [23:0]   shift_reg_426_re;
  reg        [23:0]   shift_reg_426_im;
  reg        [23:0]   shift_reg_427_re;
  reg        [23:0]   shift_reg_427_im;
  reg        [23:0]   shift_reg_428_re;
  reg        [23:0]   shift_reg_428_im;
  reg        [23:0]   shift_reg_429_re;
  reg        [23:0]   shift_reg_429_im;
  reg        [23:0]   shift_reg_430_re;
  reg        [23:0]   shift_reg_430_im;
  reg        [23:0]   shift_reg_431_re;
  reg        [23:0]   shift_reg_431_im;
  reg        [23:0]   shift_reg_432_re;
  reg        [23:0]   shift_reg_432_im;
  reg        [23:0]   shift_reg_433_re;
  reg        [23:0]   shift_reg_433_im;
  reg        [23:0]   shift_reg_434_re;
  reg        [23:0]   shift_reg_434_im;
  reg        [23:0]   shift_reg_435_re;
  reg        [23:0]   shift_reg_435_im;
  reg        [23:0]   shift_reg_436_re;
  reg        [23:0]   shift_reg_436_im;
  reg        [23:0]   shift_reg_437_re;
  reg        [23:0]   shift_reg_437_im;
  reg        [23:0]   shift_reg_438_re;
  reg        [23:0]   shift_reg_438_im;
  reg        [23:0]   shift_reg_439_re;
  reg        [23:0]   shift_reg_439_im;
  reg        [23:0]   shift_reg_440_re;
  reg        [23:0]   shift_reg_440_im;
  reg        [23:0]   shift_reg_441_re;
  reg        [23:0]   shift_reg_441_im;
  reg        [23:0]   shift_reg_442_re;
  reg        [23:0]   shift_reg_442_im;
  reg        [23:0]   shift_reg_443_re;
  reg        [23:0]   shift_reg_443_im;
  reg        [23:0]   shift_reg_444_re;
  reg        [23:0]   shift_reg_444_im;
  reg        [23:0]   shift_reg_445_re;
  reg        [23:0]   shift_reg_445_im;
  reg        [23:0]   shift_reg_446_re;
  reg        [23:0]   shift_reg_446_im;
  reg        [23:0]   shift_reg_447_re;
  reg        [23:0]   shift_reg_447_im;
  reg        [23:0]   shift_reg_448_re;
  reg        [23:0]   shift_reg_448_im;
  reg        [23:0]   shift_reg_449_re;
  reg        [23:0]   shift_reg_449_im;
  reg        [23:0]   shift_reg_450_re;
  reg        [23:0]   shift_reg_450_im;
  reg        [23:0]   shift_reg_451_re;
  reg        [23:0]   shift_reg_451_im;
  reg        [23:0]   shift_reg_452_re;
  reg        [23:0]   shift_reg_452_im;
  reg        [23:0]   shift_reg_453_re;
  reg        [23:0]   shift_reg_453_im;
  reg        [23:0]   shift_reg_454_re;
  reg        [23:0]   shift_reg_454_im;
  reg        [23:0]   shift_reg_455_re;
  reg        [23:0]   shift_reg_455_im;
  reg        [23:0]   shift_reg_456_re;
  reg        [23:0]   shift_reg_456_im;
  reg        [23:0]   shift_reg_457_re;
  reg        [23:0]   shift_reg_457_im;
  reg        [23:0]   shift_reg_458_re;
  reg        [23:0]   shift_reg_458_im;
  reg        [23:0]   shift_reg_459_re;
  reg        [23:0]   shift_reg_459_im;
  reg        [23:0]   shift_reg_460_re;
  reg        [23:0]   shift_reg_460_im;
  reg        [23:0]   shift_reg_461_re;
  reg        [23:0]   shift_reg_461_im;
  reg        [23:0]   shift_reg_462_re;
  reg        [23:0]   shift_reg_462_im;
  reg        [23:0]   shift_reg_463_re;
  reg        [23:0]   shift_reg_463_im;
  reg        [23:0]   shift_reg_464_re;
  reg        [23:0]   shift_reg_464_im;
  reg        [23:0]   shift_reg_465_re;
  reg        [23:0]   shift_reg_465_im;
  reg        [23:0]   shift_reg_466_re;
  reg        [23:0]   shift_reg_466_im;
  reg        [23:0]   shift_reg_467_re;
  reg        [23:0]   shift_reg_467_im;
  reg        [23:0]   shift_reg_468_re;
  reg        [23:0]   shift_reg_468_im;
  reg        [23:0]   shift_reg_469_re;
  reg        [23:0]   shift_reg_469_im;
  reg        [23:0]   shift_reg_470_re;
  reg        [23:0]   shift_reg_470_im;
  reg        [23:0]   shift_reg_471_re;
  reg        [23:0]   shift_reg_471_im;
  reg        [23:0]   shift_reg_472_re;
  reg        [23:0]   shift_reg_472_im;
  reg        [23:0]   shift_reg_473_re;
  reg        [23:0]   shift_reg_473_im;
  reg        [23:0]   shift_reg_474_re;
  reg        [23:0]   shift_reg_474_im;
  reg        [23:0]   shift_reg_475_re;
  reg        [23:0]   shift_reg_475_im;
  reg        [23:0]   shift_reg_476_re;
  reg        [23:0]   shift_reg_476_im;
  reg        [23:0]   shift_reg_477_re;
  reg        [23:0]   shift_reg_477_im;
  reg        [23:0]   shift_reg_478_re;
  reg        [23:0]   shift_reg_478_im;
  reg        [23:0]   shift_reg_479_re;
  reg        [23:0]   shift_reg_479_im;
  reg        [23:0]   shift_reg_480_re;
  reg        [23:0]   shift_reg_480_im;
  reg        [23:0]   shift_reg_481_re;
  reg        [23:0]   shift_reg_481_im;
  reg        [23:0]   shift_reg_482_re;
  reg        [23:0]   shift_reg_482_im;
  reg        [23:0]   shift_reg_483_re;
  reg        [23:0]   shift_reg_483_im;
  reg        [23:0]   shift_reg_484_re;
  reg        [23:0]   shift_reg_484_im;
  reg        [23:0]   shift_reg_485_re;
  reg        [23:0]   shift_reg_485_im;
  reg        [23:0]   shift_reg_486_re;
  reg        [23:0]   shift_reg_486_im;
  reg        [23:0]   shift_reg_487_re;
  reg        [23:0]   shift_reg_487_im;
  reg        [23:0]   shift_reg_488_re;
  reg        [23:0]   shift_reg_488_im;
  reg        [23:0]   shift_reg_489_re;
  reg        [23:0]   shift_reg_489_im;
  reg        [23:0]   shift_reg_490_re;
  reg        [23:0]   shift_reg_490_im;
  reg        [23:0]   shift_reg_491_re;
  reg        [23:0]   shift_reg_491_im;
  reg        [23:0]   shift_reg_492_re;
  reg        [23:0]   shift_reg_492_im;
  reg        [23:0]   shift_reg_493_re;
  reg        [23:0]   shift_reg_493_im;
  reg        [23:0]   shift_reg_494_re;
  reg        [23:0]   shift_reg_494_im;
  reg        [23:0]   shift_reg_495_re;
  reg        [23:0]   shift_reg_495_im;
  reg        [23:0]   shift_reg_496_re;
  reg        [23:0]   shift_reg_496_im;
  reg        [23:0]   shift_reg_497_re;
  reg        [23:0]   shift_reg_497_im;
  reg        [23:0]   shift_reg_498_re;
  reg        [23:0]   shift_reg_498_im;
  reg        [23:0]   shift_reg_499_re;
  reg        [23:0]   shift_reg_499_im;
  reg        [23:0]   shift_reg_500_re;
  reg        [23:0]   shift_reg_500_im;
  reg        [23:0]   shift_reg_501_re;
  reg        [23:0]   shift_reg_501_im;
  reg        [23:0]   shift_reg_502_re;
  reg        [23:0]   shift_reg_502_im;
  reg        [23:0]   shift_reg_503_re;
  reg        [23:0]   shift_reg_503_im;
  reg        [23:0]   shift_reg_504_re;
  reg        [23:0]   shift_reg_504_im;
  reg        [23:0]   shift_reg_505_re;
  reg        [23:0]   shift_reg_505_im;
  reg        [23:0]   shift_reg_506_re;
  reg        [23:0]   shift_reg_506_im;
  reg        [23:0]   shift_reg_507_re;
  reg        [23:0]   shift_reg_507_im;
  reg        [23:0]   shift_reg_508_re;
  reg        [23:0]   shift_reg_508_im;
  reg        [23:0]   shift_reg_509_re;
  reg        [23:0]   shift_reg_509_im;
  reg        [23:0]   shift_reg_510_re;
  reg        [23:0]   shift_reg_510_im;
  reg        [23:0]   shift_reg_511_re;
  reg        [23:0]   shift_reg_511_im;
  reg        [23:0]   shift_reg_512_re;
  reg        [23:0]   shift_reg_512_im;
  reg        [23:0]   shift_reg_513_re;
  reg        [23:0]   shift_reg_513_im;
  reg        [23:0]   shift_reg_514_re;
  reg        [23:0]   shift_reg_514_im;
  reg        [23:0]   shift_reg_515_re;
  reg        [23:0]   shift_reg_515_im;
  reg        [23:0]   shift_reg_516_re;
  reg        [23:0]   shift_reg_516_im;
  reg        [23:0]   shift_reg_517_re;
  reg        [23:0]   shift_reg_517_im;
  reg        [23:0]   shift_reg_518_re;
  reg        [23:0]   shift_reg_518_im;
  reg        [23:0]   shift_reg_519_re;
  reg        [23:0]   shift_reg_519_im;
  reg        [23:0]   shift_reg_520_re;
  reg        [23:0]   shift_reg_520_im;
  reg        [23:0]   shift_reg_521_re;
  reg        [23:0]   shift_reg_521_im;
  reg        [23:0]   shift_reg_522_re;
  reg        [23:0]   shift_reg_522_im;
  reg        [23:0]   shift_reg_523_re;
  reg        [23:0]   shift_reg_523_im;
  reg        [23:0]   shift_reg_524_re;
  reg        [23:0]   shift_reg_524_im;
  reg        [23:0]   shift_reg_525_re;
  reg        [23:0]   shift_reg_525_im;
  reg        [23:0]   shift_reg_526_re;
  reg        [23:0]   shift_reg_526_im;
  reg        [23:0]   shift_reg_527_re;
  reg        [23:0]   shift_reg_527_im;
  reg        [23:0]   shift_reg_528_re;
  reg        [23:0]   shift_reg_528_im;
  reg        [23:0]   shift_reg_529_re;
  reg        [23:0]   shift_reg_529_im;
  reg        [23:0]   shift_reg_530_re;
  reg        [23:0]   shift_reg_530_im;
  reg        [23:0]   shift_reg_531_re;
  reg        [23:0]   shift_reg_531_im;
  reg        [23:0]   shift_reg_532_re;
  reg        [23:0]   shift_reg_532_im;
  reg        [23:0]   shift_reg_533_re;
  reg        [23:0]   shift_reg_533_im;
  reg        [23:0]   shift_reg_534_re;
  reg        [23:0]   shift_reg_534_im;
  reg        [23:0]   shift_reg_535_re;
  reg        [23:0]   shift_reg_535_im;
  reg        [23:0]   shift_reg_536_re;
  reg        [23:0]   shift_reg_536_im;
  reg        [23:0]   shift_reg_537_re;
  reg        [23:0]   shift_reg_537_im;
  reg        [23:0]   shift_reg_538_re;
  reg        [23:0]   shift_reg_538_im;
  reg        [23:0]   shift_reg_539_re;
  reg        [23:0]   shift_reg_539_im;
  reg        [23:0]   shift_reg_540_re;
  reg        [23:0]   shift_reg_540_im;
  reg        [23:0]   shift_reg_541_re;
  reg        [23:0]   shift_reg_541_im;
  reg        [23:0]   shift_reg_542_re;
  reg        [23:0]   shift_reg_542_im;
  reg        [23:0]   shift_reg_543_re;
  reg        [23:0]   shift_reg_543_im;
  reg        [23:0]   shift_reg_544_re;
  reg        [23:0]   shift_reg_544_im;
  reg        [23:0]   shift_reg_545_re;
  reg        [23:0]   shift_reg_545_im;
  reg        [23:0]   shift_reg_546_re;
  reg        [23:0]   shift_reg_546_im;
  reg        [23:0]   shift_reg_547_re;
  reg        [23:0]   shift_reg_547_im;
  reg        [23:0]   shift_reg_548_re;
  reg        [23:0]   shift_reg_548_im;
  reg        [23:0]   shift_reg_549_re;
  reg        [23:0]   shift_reg_549_im;
  reg        [23:0]   shift_reg_550_re;
  reg        [23:0]   shift_reg_550_im;
  reg        [23:0]   shift_reg_551_re;
  reg        [23:0]   shift_reg_551_im;
  reg        [23:0]   shift_reg_552_re;
  reg        [23:0]   shift_reg_552_im;
  reg        [23:0]   shift_reg_553_re;
  reg        [23:0]   shift_reg_553_im;
  reg        [23:0]   shift_reg_554_re;
  reg        [23:0]   shift_reg_554_im;
  reg        [23:0]   shift_reg_555_re;
  reg        [23:0]   shift_reg_555_im;
  reg        [23:0]   shift_reg_556_re;
  reg        [23:0]   shift_reg_556_im;
  reg        [23:0]   shift_reg_557_re;
  reg        [23:0]   shift_reg_557_im;
  reg        [23:0]   shift_reg_558_re;
  reg        [23:0]   shift_reg_558_im;
  reg        [23:0]   shift_reg_559_re;
  reg        [23:0]   shift_reg_559_im;
  reg        [23:0]   shift_reg_560_re;
  reg        [23:0]   shift_reg_560_im;
  reg        [23:0]   shift_reg_561_re;
  reg        [23:0]   shift_reg_561_im;
  reg        [23:0]   shift_reg_562_re;
  reg        [23:0]   shift_reg_562_im;
  reg        [23:0]   shift_reg_563_re;
  reg        [23:0]   shift_reg_563_im;
  reg        [23:0]   shift_reg_564_re;
  reg        [23:0]   shift_reg_564_im;
  reg        [23:0]   shift_reg_565_re;
  reg        [23:0]   shift_reg_565_im;
  reg        [23:0]   shift_reg_566_re;
  reg        [23:0]   shift_reg_566_im;
  reg        [23:0]   shift_reg_567_re;
  reg        [23:0]   shift_reg_567_im;
  reg        [23:0]   shift_reg_568_re;
  reg        [23:0]   shift_reg_568_im;
  reg        [23:0]   shift_reg_569_re;
  reg        [23:0]   shift_reg_569_im;
  reg        [23:0]   shift_reg_570_re;
  reg        [23:0]   shift_reg_570_im;
  reg        [23:0]   shift_reg_571_re;
  reg        [23:0]   shift_reg_571_im;
  reg        [23:0]   shift_reg_572_re;
  reg        [23:0]   shift_reg_572_im;
  reg        [23:0]   shift_reg_573_re;
  reg        [23:0]   shift_reg_573_im;
  reg        [23:0]   shift_reg_574_re;
  reg        [23:0]   shift_reg_574_im;
  reg        [23:0]   shift_reg_575_re;
  reg        [23:0]   shift_reg_575_im;
  reg        [23:0]   shift_reg_576_re;
  reg        [23:0]   shift_reg_576_im;
  reg        [23:0]   shift_reg_577_re;
  reg        [23:0]   shift_reg_577_im;
  reg        [23:0]   shift_reg_578_re;
  reg        [23:0]   shift_reg_578_im;
  reg        [23:0]   shift_reg_579_re;
  reg        [23:0]   shift_reg_579_im;
  reg        [23:0]   shift_reg_580_re;
  reg        [23:0]   shift_reg_580_im;
  reg        [23:0]   shift_reg_581_re;
  reg        [23:0]   shift_reg_581_im;
  reg        [23:0]   shift_reg_582_re;
  reg        [23:0]   shift_reg_582_im;
  reg        [23:0]   shift_reg_583_re;
  reg        [23:0]   shift_reg_583_im;
  reg        [23:0]   shift_reg_584_re;
  reg        [23:0]   shift_reg_584_im;
  reg        [23:0]   shift_reg_585_re;
  reg        [23:0]   shift_reg_585_im;
  reg        [23:0]   shift_reg_586_re;
  reg        [23:0]   shift_reg_586_im;
  reg        [23:0]   shift_reg_587_re;
  reg        [23:0]   shift_reg_587_im;
  reg        [23:0]   shift_reg_588_re;
  reg        [23:0]   shift_reg_588_im;
  reg        [23:0]   shift_reg_589_re;
  reg        [23:0]   shift_reg_589_im;
  reg        [23:0]   shift_reg_590_re;
  reg        [23:0]   shift_reg_590_im;
  reg        [23:0]   shift_reg_591_re;
  reg        [23:0]   shift_reg_591_im;
  reg        [23:0]   shift_reg_592_re;
  reg        [23:0]   shift_reg_592_im;
  reg        [23:0]   shift_reg_593_re;
  reg        [23:0]   shift_reg_593_im;
  reg        [23:0]   shift_reg_594_re;
  reg        [23:0]   shift_reg_594_im;
  reg        [23:0]   shift_reg_595_re;
  reg        [23:0]   shift_reg_595_im;
  reg        [23:0]   shift_reg_596_re;
  reg        [23:0]   shift_reg_596_im;
  reg        [23:0]   shift_reg_597_re;
  reg        [23:0]   shift_reg_597_im;
  reg        [23:0]   shift_reg_598_re;
  reg        [23:0]   shift_reg_598_im;
  reg        [23:0]   shift_reg_599_re;
  reg        [23:0]   shift_reg_599_im;
  reg        [23:0]   shift_reg_600_re;
  reg        [23:0]   shift_reg_600_im;
  reg        [23:0]   shift_reg_601_re;
  reg        [23:0]   shift_reg_601_im;
  reg        [23:0]   shift_reg_602_re;
  reg        [23:0]   shift_reg_602_im;
  reg        [23:0]   shift_reg_603_re;
  reg        [23:0]   shift_reg_603_im;
  reg        [23:0]   shift_reg_604_re;
  reg        [23:0]   shift_reg_604_im;
  reg        [23:0]   shift_reg_605_re;
  reg        [23:0]   shift_reg_605_im;
  reg        [23:0]   shift_reg_606_re;
  reg        [23:0]   shift_reg_606_im;
  reg        [23:0]   shift_reg_607_re;
  reg        [23:0]   shift_reg_607_im;
  reg        [23:0]   shift_reg_608_re;
  reg        [23:0]   shift_reg_608_im;
  reg        [23:0]   shift_reg_609_re;
  reg        [23:0]   shift_reg_609_im;
  reg        [23:0]   shift_reg_610_re;
  reg        [23:0]   shift_reg_610_im;
  reg        [23:0]   shift_reg_611_re;
  reg        [23:0]   shift_reg_611_im;
  reg        [23:0]   shift_reg_612_re;
  reg        [23:0]   shift_reg_612_im;
  reg        [23:0]   shift_reg_613_re;
  reg        [23:0]   shift_reg_613_im;
  reg        [23:0]   shift_reg_614_re;
  reg        [23:0]   shift_reg_614_im;
  reg        [23:0]   shift_reg_615_re;
  reg        [23:0]   shift_reg_615_im;
  reg        [23:0]   shift_reg_616_re;
  reg        [23:0]   shift_reg_616_im;
  reg        [23:0]   shift_reg_617_re;
  reg        [23:0]   shift_reg_617_im;
  reg        [23:0]   shift_reg_618_re;
  reg        [23:0]   shift_reg_618_im;
  reg        [23:0]   shift_reg_619_re;
  reg        [23:0]   shift_reg_619_im;
  reg        [23:0]   shift_reg_620_re;
  reg        [23:0]   shift_reg_620_im;
  reg        [23:0]   shift_reg_621_re;
  reg        [23:0]   shift_reg_621_im;
  reg        [23:0]   shift_reg_622_re;
  reg        [23:0]   shift_reg_622_im;
  reg        [23:0]   shift_reg_623_re;
  reg        [23:0]   shift_reg_623_im;
  reg        [23:0]   shift_reg_624_re;
  reg        [23:0]   shift_reg_624_im;
  reg        [23:0]   shift_reg_625_re;
  reg        [23:0]   shift_reg_625_im;
  reg        [23:0]   shift_reg_626_re;
  reg        [23:0]   shift_reg_626_im;
  reg        [23:0]   shift_reg_627_re;
  reg        [23:0]   shift_reg_627_im;
  reg        [23:0]   shift_reg_628_re;
  reg        [23:0]   shift_reg_628_im;
  reg        [23:0]   shift_reg_629_re;
  reg        [23:0]   shift_reg_629_im;
  reg        [23:0]   shift_reg_630_re;
  reg        [23:0]   shift_reg_630_im;
  reg        [23:0]   shift_reg_631_re;
  reg        [23:0]   shift_reg_631_im;
  reg        [23:0]   shift_reg_632_re;
  reg        [23:0]   shift_reg_632_im;
  reg        [23:0]   shift_reg_633_re;
  reg        [23:0]   shift_reg_633_im;
  reg        [23:0]   shift_reg_634_re;
  reg        [23:0]   shift_reg_634_im;
  reg        [23:0]   shift_reg_635_re;
  reg        [23:0]   shift_reg_635_im;
  reg        [23:0]   shift_reg_636_re;
  reg        [23:0]   shift_reg_636_im;
  reg        [23:0]   shift_reg_637_re;
  reg        [23:0]   shift_reg_637_im;
  reg        [23:0]   shift_reg_638_re;
  reg        [23:0]   shift_reg_638_im;
  reg        [23:0]   shift_reg_639_re;
  reg        [23:0]   shift_reg_639_im;
  reg        [23:0]   shift_reg_640_re;
  reg        [23:0]   shift_reg_640_im;
  reg        [23:0]   shift_reg_641_re;
  reg        [23:0]   shift_reg_641_im;
  reg        [23:0]   shift_reg_642_re;
  reg        [23:0]   shift_reg_642_im;
  reg        [23:0]   shift_reg_643_re;
  reg        [23:0]   shift_reg_643_im;
  reg        [23:0]   shift_reg_644_re;
  reg        [23:0]   shift_reg_644_im;
  reg        [23:0]   shift_reg_645_re;
  reg        [23:0]   shift_reg_645_im;
  reg        [23:0]   shift_reg_646_re;
  reg        [23:0]   shift_reg_646_im;
  reg        [23:0]   shift_reg_647_re;
  reg        [23:0]   shift_reg_647_im;
  reg        [23:0]   shift_reg_648_re;
  reg        [23:0]   shift_reg_648_im;
  reg        [23:0]   shift_reg_649_re;
  reg        [23:0]   shift_reg_649_im;
  reg        [23:0]   shift_reg_650_re;
  reg        [23:0]   shift_reg_650_im;
  reg        [23:0]   shift_reg_651_re;
  reg        [23:0]   shift_reg_651_im;
  reg        [23:0]   shift_reg_652_re;
  reg        [23:0]   shift_reg_652_im;
  reg        [23:0]   shift_reg_653_re;
  reg        [23:0]   shift_reg_653_im;
  reg        [23:0]   shift_reg_654_re;
  reg        [23:0]   shift_reg_654_im;
  reg        [23:0]   shift_reg_655_re;
  reg        [23:0]   shift_reg_655_im;
  reg        [23:0]   shift_reg_656_re;
  reg        [23:0]   shift_reg_656_im;
  reg        [23:0]   shift_reg_657_re;
  reg        [23:0]   shift_reg_657_im;
  reg        [23:0]   shift_reg_658_re;
  reg        [23:0]   shift_reg_658_im;
  reg        [23:0]   shift_reg_659_re;
  reg        [23:0]   shift_reg_659_im;
  reg        [23:0]   shift_reg_660_re;
  reg        [23:0]   shift_reg_660_im;
  reg        [23:0]   shift_reg_661_re;
  reg        [23:0]   shift_reg_661_im;
  reg        [23:0]   shift_reg_662_re;
  reg        [23:0]   shift_reg_662_im;
  reg        [23:0]   shift_reg_663_re;
  reg        [23:0]   shift_reg_663_im;
  reg        [23:0]   shift_reg_664_re;
  reg        [23:0]   shift_reg_664_im;
  reg        [23:0]   shift_reg_665_re;
  reg        [23:0]   shift_reg_665_im;
  reg        [23:0]   shift_reg_666_re;
  reg        [23:0]   shift_reg_666_im;
  reg        [23:0]   shift_reg_667_re;
  reg        [23:0]   shift_reg_667_im;
  reg        [23:0]   shift_reg_668_re;
  reg        [23:0]   shift_reg_668_im;
  reg        [23:0]   shift_reg_669_re;
  reg        [23:0]   shift_reg_669_im;
  reg        [23:0]   shift_reg_670_re;
  reg        [23:0]   shift_reg_670_im;
  reg        [23:0]   shift_reg_671_re;
  reg        [23:0]   shift_reg_671_im;
  reg        [23:0]   shift_reg_672_re;
  reg        [23:0]   shift_reg_672_im;
  reg        [23:0]   shift_reg_673_re;
  reg        [23:0]   shift_reg_673_im;
  reg        [23:0]   shift_reg_674_re;
  reg        [23:0]   shift_reg_674_im;
  reg        [23:0]   shift_reg_675_re;
  reg        [23:0]   shift_reg_675_im;
  reg        [23:0]   shift_reg_676_re;
  reg        [23:0]   shift_reg_676_im;
  reg        [23:0]   shift_reg_677_re;
  reg        [23:0]   shift_reg_677_im;
  reg        [23:0]   shift_reg_678_re;
  reg        [23:0]   shift_reg_678_im;
  reg        [23:0]   shift_reg_679_re;
  reg        [23:0]   shift_reg_679_im;
  reg        [23:0]   shift_reg_680_re;
  reg        [23:0]   shift_reg_680_im;
  reg        [23:0]   shift_reg_681_re;
  reg        [23:0]   shift_reg_681_im;
  reg        [23:0]   shift_reg_682_re;
  reg        [23:0]   shift_reg_682_im;
  reg        [23:0]   shift_reg_683_re;
  reg        [23:0]   shift_reg_683_im;
  reg        [23:0]   shift_reg_684_re;
  reg        [23:0]   shift_reg_684_im;
  reg        [23:0]   shift_reg_685_re;
  reg        [23:0]   shift_reg_685_im;
  reg        [23:0]   shift_reg_686_re;
  reg        [23:0]   shift_reg_686_im;
  reg        [23:0]   shift_reg_687_re;
  reg        [23:0]   shift_reg_687_im;
  reg        [23:0]   shift_reg_688_re;
  reg        [23:0]   shift_reg_688_im;
  reg        [23:0]   shift_reg_689_re;
  reg        [23:0]   shift_reg_689_im;
  reg        [23:0]   shift_reg_690_re;
  reg        [23:0]   shift_reg_690_im;
  reg        [23:0]   shift_reg_691_re;
  reg        [23:0]   shift_reg_691_im;
  reg        [23:0]   shift_reg_692_re;
  reg        [23:0]   shift_reg_692_im;
  reg        [23:0]   shift_reg_693_re;
  reg        [23:0]   shift_reg_693_im;
  reg        [23:0]   shift_reg_694_re;
  reg        [23:0]   shift_reg_694_im;
  reg        [23:0]   shift_reg_695_re;
  reg        [23:0]   shift_reg_695_im;
  reg        [23:0]   shift_reg_696_re;
  reg        [23:0]   shift_reg_696_im;
  reg        [23:0]   shift_reg_697_re;
  reg        [23:0]   shift_reg_697_im;
  reg        [23:0]   shift_reg_698_re;
  reg        [23:0]   shift_reg_698_im;
  reg        [23:0]   shift_reg_699_re;
  reg        [23:0]   shift_reg_699_im;
  reg        [23:0]   shift_reg_700_re;
  reg        [23:0]   shift_reg_700_im;
  reg        [23:0]   shift_reg_701_re;
  reg        [23:0]   shift_reg_701_im;
  reg        [23:0]   shift_reg_702_re;
  reg        [23:0]   shift_reg_702_im;
  reg        [23:0]   shift_reg_703_re;
  reg        [23:0]   shift_reg_703_im;
  reg        [23:0]   shift_reg_704_re;
  reg        [23:0]   shift_reg_704_im;
  reg        [23:0]   shift_reg_705_re;
  reg        [23:0]   shift_reg_705_im;
  reg        [23:0]   shift_reg_706_re;
  reg        [23:0]   shift_reg_706_im;
  reg        [23:0]   shift_reg_707_re;
  reg        [23:0]   shift_reg_707_im;
  reg        [23:0]   shift_reg_708_re;
  reg        [23:0]   shift_reg_708_im;
  reg        [23:0]   shift_reg_709_re;
  reg        [23:0]   shift_reg_709_im;
  reg        [23:0]   shift_reg_710_re;
  reg        [23:0]   shift_reg_710_im;
  reg        [23:0]   shift_reg_711_re;
  reg        [23:0]   shift_reg_711_im;
  reg        [23:0]   shift_reg_712_re;
  reg        [23:0]   shift_reg_712_im;
  reg        [23:0]   shift_reg_713_re;
  reg        [23:0]   shift_reg_713_im;
  reg        [23:0]   shift_reg_714_re;
  reg        [23:0]   shift_reg_714_im;
  reg        [23:0]   shift_reg_715_re;
  reg        [23:0]   shift_reg_715_im;
  reg        [23:0]   shift_reg_716_re;
  reg        [23:0]   shift_reg_716_im;
  reg        [23:0]   shift_reg_717_re;
  reg        [23:0]   shift_reg_717_im;
  reg        [23:0]   shift_reg_718_re;
  reg        [23:0]   shift_reg_718_im;
  reg        [23:0]   shift_reg_719_re;
  reg        [23:0]   shift_reg_719_im;
  reg        [23:0]   shift_reg_720_re;
  reg        [23:0]   shift_reg_720_im;
  reg        [23:0]   shift_reg_721_re;
  reg        [23:0]   shift_reg_721_im;
  reg        [23:0]   shift_reg_722_re;
  reg        [23:0]   shift_reg_722_im;
  reg        [23:0]   shift_reg_723_re;
  reg        [23:0]   shift_reg_723_im;
  reg        [23:0]   shift_reg_724_re;
  reg        [23:0]   shift_reg_724_im;
  reg        [23:0]   shift_reg_725_re;
  reg        [23:0]   shift_reg_725_im;
  reg        [23:0]   shift_reg_726_re;
  reg        [23:0]   shift_reg_726_im;
  reg        [23:0]   shift_reg_727_re;
  reg        [23:0]   shift_reg_727_im;
  reg        [23:0]   shift_reg_728_re;
  reg        [23:0]   shift_reg_728_im;
  reg        [23:0]   shift_reg_729_re;
  reg        [23:0]   shift_reg_729_im;
  reg        [23:0]   shift_reg_730_re;
  reg        [23:0]   shift_reg_730_im;
  reg        [23:0]   shift_reg_731_re;
  reg        [23:0]   shift_reg_731_im;
  reg        [23:0]   shift_reg_732_re;
  reg        [23:0]   shift_reg_732_im;
  reg        [23:0]   shift_reg_733_re;
  reg        [23:0]   shift_reg_733_im;
  reg        [23:0]   shift_reg_734_re;
  reg        [23:0]   shift_reg_734_im;
  reg        [23:0]   shift_reg_735_re;
  reg        [23:0]   shift_reg_735_im;
  reg        [23:0]   shift_reg_736_re;
  reg        [23:0]   shift_reg_736_im;
  reg        [23:0]   shift_reg_737_re;
  reg        [23:0]   shift_reg_737_im;
  reg        [23:0]   shift_reg_738_re;
  reg        [23:0]   shift_reg_738_im;
  reg        [23:0]   shift_reg_739_re;
  reg        [23:0]   shift_reg_739_im;
  reg        [23:0]   shift_reg_740_re;
  reg        [23:0]   shift_reg_740_im;
  reg        [23:0]   shift_reg_741_re;
  reg        [23:0]   shift_reg_741_im;
  reg        [23:0]   shift_reg_742_re;
  reg        [23:0]   shift_reg_742_im;
  reg        [23:0]   shift_reg_743_re;
  reg        [23:0]   shift_reg_743_im;
  reg        [23:0]   shift_reg_744_re;
  reg        [23:0]   shift_reg_744_im;
  reg        [23:0]   shift_reg_745_re;
  reg        [23:0]   shift_reg_745_im;
  reg        [23:0]   shift_reg_746_re;
  reg        [23:0]   shift_reg_746_im;
  reg        [23:0]   shift_reg_747_re;
  reg        [23:0]   shift_reg_747_im;
  reg        [23:0]   shift_reg_748_re;
  reg        [23:0]   shift_reg_748_im;
  reg        [23:0]   shift_reg_749_re;
  reg        [23:0]   shift_reg_749_im;
  reg        [23:0]   shift_reg_750_re;
  reg        [23:0]   shift_reg_750_im;
  reg        [23:0]   shift_reg_751_re;
  reg        [23:0]   shift_reg_751_im;
  reg        [23:0]   shift_reg_752_re;
  reg        [23:0]   shift_reg_752_im;
  reg        [23:0]   shift_reg_753_re;
  reg        [23:0]   shift_reg_753_im;
  reg        [23:0]   shift_reg_754_re;
  reg        [23:0]   shift_reg_754_im;
  reg        [23:0]   shift_reg_755_re;
  reg        [23:0]   shift_reg_755_im;
  reg        [23:0]   shift_reg_756_re;
  reg        [23:0]   shift_reg_756_im;
  reg        [23:0]   shift_reg_757_re;
  reg        [23:0]   shift_reg_757_im;
  reg        [23:0]   shift_reg_758_re;
  reg        [23:0]   shift_reg_758_im;
  reg        [23:0]   shift_reg_759_re;
  reg        [23:0]   shift_reg_759_im;
  reg        [23:0]   shift_reg_760_re;
  reg        [23:0]   shift_reg_760_im;
  reg        [23:0]   shift_reg_761_re;
  reg        [23:0]   shift_reg_761_im;
  reg        [23:0]   shift_reg_762_re;
  reg        [23:0]   shift_reg_762_im;
  reg        [23:0]   shift_reg_763_re;
  reg        [23:0]   shift_reg_763_im;
  reg        [23:0]   shift_reg_764_re;
  reg        [23:0]   shift_reg_764_im;
  reg        [23:0]   shift_reg_765_re;
  reg        [23:0]   shift_reg_765_im;
  reg        [23:0]   shift_reg_766_re;
  reg        [23:0]   shift_reg_766_im;
  reg        [23:0]   shift_reg_767_re;
  reg        [23:0]   shift_reg_767_im;
  reg        [23:0]   shift_reg_768_re;
  reg        [23:0]   shift_reg_768_im;
  reg        [23:0]   shift_reg_769_re;
  reg        [23:0]   shift_reg_769_im;
  reg        [23:0]   shift_reg_770_re;
  reg        [23:0]   shift_reg_770_im;
  reg        [23:0]   shift_reg_771_re;
  reg        [23:0]   shift_reg_771_im;
  reg        [23:0]   shift_reg_772_re;
  reg        [23:0]   shift_reg_772_im;
  reg        [23:0]   shift_reg_773_re;
  reg        [23:0]   shift_reg_773_im;
  reg        [23:0]   shift_reg_774_re;
  reg        [23:0]   shift_reg_774_im;
  reg        [23:0]   shift_reg_775_re;
  reg        [23:0]   shift_reg_775_im;
  reg        [23:0]   shift_reg_776_re;
  reg        [23:0]   shift_reg_776_im;
  reg        [23:0]   shift_reg_777_re;
  reg        [23:0]   shift_reg_777_im;
  reg        [23:0]   shift_reg_778_re;
  reg        [23:0]   shift_reg_778_im;
  reg        [23:0]   shift_reg_779_re;
  reg        [23:0]   shift_reg_779_im;
  reg        [23:0]   shift_reg_780_re;
  reg        [23:0]   shift_reg_780_im;
  reg        [23:0]   shift_reg_781_re;
  reg        [23:0]   shift_reg_781_im;
  reg        [23:0]   shift_reg_782_re;
  reg        [23:0]   shift_reg_782_im;
  reg        [23:0]   shift_reg_783_re;
  reg        [23:0]   shift_reg_783_im;
  reg        [23:0]   shift_reg_784_re;
  reg        [23:0]   shift_reg_784_im;
  reg        [23:0]   shift_reg_785_re;
  reg        [23:0]   shift_reg_785_im;
  reg        [23:0]   shift_reg_786_re;
  reg        [23:0]   shift_reg_786_im;
  reg        [23:0]   shift_reg_787_re;
  reg        [23:0]   shift_reg_787_im;
  reg        [23:0]   shift_reg_788_re;
  reg        [23:0]   shift_reg_788_im;
  reg        [23:0]   shift_reg_789_re;
  reg        [23:0]   shift_reg_789_im;
  reg        [23:0]   shift_reg_790_re;
  reg        [23:0]   shift_reg_790_im;
  reg        [23:0]   shift_reg_791_re;
  reg        [23:0]   shift_reg_791_im;
  reg        [23:0]   shift_reg_792_re;
  reg        [23:0]   shift_reg_792_im;
  reg        [23:0]   shift_reg_793_re;
  reg        [23:0]   shift_reg_793_im;
  reg        [23:0]   shift_reg_794_re;
  reg        [23:0]   shift_reg_794_im;
  reg        [23:0]   shift_reg_795_re;
  reg        [23:0]   shift_reg_795_im;
  reg        [23:0]   shift_reg_796_re;
  reg        [23:0]   shift_reg_796_im;
  reg        [23:0]   shift_reg_797_re;
  reg        [23:0]   shift_reg_797_im;
  reg        [23:0]   shift_reg_798_re;
  reg        [23:0]   shift_reg_798_im;
  reg        [23:0]   shift_reg_799_re;
  reg        [23:0]   shift_reg_799_im;
  reg        [23:0]   shift_reg_800_re;
  reg        [23:0]   shift_reg_800_im;
  reg        [23:0]   shift_reg_801_re;
  reg        [23:0]   shift_reg_801_im;
  reg        [23:0]   shift_reg_802_re;
  reg        [23:0]   shift_reg_802_im;
  reg        [23:0]   shift_reg_803_re;
  reg        [23:0]   shift_reg_803_im;
  reg        [23:0]   shift_reg_804_re;
  reg        [23:0]   shift_reg_804_im;
  reg        [23:0]   shift_reg_805_re;
  reg        [23:0]   shift_reg_805_im;
  reg        [23:0]   shift_reg_806_re;
  reg        [23:0]   shift_reg_806_im;
  reg        [23:0]   shift_reg_807_re;
  reg        [23:0]   shift_reg_807_im;
  reg        [23:0]   shift_reg_808_re;
  reg        [23:0]   shift_reg_808_im;
  reg        [23:0]   shift_reg_809_re;
  reg        [23:0]   shift_reg_809_im;
  reg        [23:0]   shift_reg_810_re;
  reg        [23:0]   shift_reg_810_im;
  reg        [23:0]   shift_reg_811_re;
  reg        [23:0]   shift_reg_811_im;
  reg        [23:0]   shift_reg_812_re;
  reg        [23:0]   shift_reg_812_im;
  reg        [23:0]   shift_reg_813_re;
  reg        [23:0]   shift_reg_813_im;
  reg        [23:0]   shift_reg_814_re;
  reg        [23:0]   shift_reg_814_im;
  reg        [23:0]   shift_reg_815_re;
  reg        [23:0]   shift_reg_815_im;
  reg        [23:0]   shift_reg_816_re;
  reg        [23:0]   shift_reg_816_im;
  reg        [23:0]   shift_reg_817_re;
  reg        [23:0]   shift_reg_817_im;
  reg        [23:0]   shift_reg_818_re;
  reg        [23:0]   shift_reg_818_im;
  reg        [23:0]   shift_reg_819_re;
  reg        [23:0]   shift_reg_819_im;
  reg        [23:0]   shift_reg_820_re;
  reg        [23:0]   shift_reg_820_im;
  reg        [23:0]   shift_reg_821_re;
  reg        [23:0]   shift_reg_821_im;
  reg        [23:0]   shift_reg_822_re;
  reg        [23:0]   shift_reg_822_im;
  reg        [23:0]   shift_reg_823_re;
  reg        [23:0]   shift_reg_823_im;
  reg        [23:0]   shift_reg_824_re;
  reg        [23:0]   shift_reg_824_im;
  reg        [23:0]   shift_reg_825_re;
  reg        [23:0]   shift_reg_825_im;
  reg        [23:0]   shift_reg_826_re;
  reg        [23:0]   shift_reg_826_im;
  reg        [23:0]   shift_reg_827_re;
  reg        [23:0]   shift_reg_827_im;
  reg        [23:0]   shift_reg_828_re;
  reg        [23:0]   shift_reg_828_im;
  reg        [23:0]   shift_reg_829_re;
  reg        [23:0]   shift_reg_829_im;
  reg        [23:0]   shift_reg_830_re;
  reg        [23:0]   shift_reg_830_im;
  reg        [23:0]   shift_reg_831_re;
  reg        [23:0]   shift_reg_831_im;
  reg        [23:0]   shift_reg_832_re;
  reg        [23:0]   shift_reg_832_im;
  reg        [23:0]   shift_reg_833_re;
  reg        [23:0]   shift_reg_833_im;
  reg        [23:0]   shift_reg_834_re;
  reg        [23:0]   shift_reg_834_im;
  reg        [23:0]   shift_reg_835_re;
  reg        [23:0]   shift_reg_835_im;
  reg        [23:0]   shift_reg_836_re;
  reg        [23:0]   shift_reg_836_im;
  reg        [23:0]   shift_reg_837_re;
  reg        [23:0]   shift_reg_837_im;
  reg        [23:0]   shift_reg_838_re;
  reg        [23:0]   shift_reg_838_im;
  reg        [23:0]   shift_reg_839_re;
  reg        [23:0]   shift_reg_839_im;
  reg        [23:0]   shift_reg_840_re;
  reg        [23:0]   shift_reg_840_im;
  reg        [23:0]   shift_reg_841_re;
  reg        [23:0]   shift_reg_841_im;
  reg        [23:0]   shift_reg_842_re;
  reg        [23:0]   shift_reg_842_im;
  reg        [23:0]   shift_reg_843_re;
  reg        [23:0]   shift_reg_843_im;
  reg        [23:0]   shift_reg_844_re;
  reg        [23:0]   shift_reg_844_im;
  reg        [23:0]   shift_reg_845_re;
  reg        [23:0]   shift_reg_845_im;
  reg        [23:0]   shift_reg_846_re;
  reg        [23:0]   shift_reg_846_im;
  reg        [23:0]   shift_reg_847_re;
  reg        [23:0]   shift_reg_847_im;
  reg        [23:0]   shift_reg_848_re;
  reg        [23:0]   shift_reg_848_im;
  reg        [23:0]   shift_reg_849_re;
  reg        [23:0]   shift_reg_849_im;
  reg        [23:0]   shift_reg_850_re;
  reg        [23:0]   shift_reg_850_im;
  reg        [23:0]   shift_reg_851_re;
  reg        [23:0]   shift_reg_851_im;
  reg        [23:0]   shift_reg_852_re;
  reg        [23:0]   shift_reg_852_im;
  reg        [23:0]   shift_reg_853_re;
  reg        [23:0]   shift_reg_853_im;
  reg        [23:0]   shift_reg_854_re;
  reg        [23:0]   shift_reg_854_im;
  reg        [23:0]   shift_reg_855_re;
  reg        [23:0]   shift_reg_855_im;
  reg        [23:0]   shift_reg_856_re;
  reg        [23:0]   shift_reg_856_im;
  reg        [23:0]   shift_reg_857_re;
  reg        [23:0]   shift_reg_857_im;
  reg        [23:0]   shift_reg_858_re;
  reg        [23:0]   shift_reg_858_im;
  reg        [23:0]   shift_reg_859_re;
  reg        [23:0]   shift_reg_859_im;
  reg        [23:0]   shift_reg_860_re;
  reg        [23:0]   shift_reg_860_im;
  reg        [23:0]   shift_reg_861_re;
  reg        [23:0]   shift_reg_861_im;
  reg        [23:0]   shift_reg_862_re;
  reg        [23:0]   shift_reg_862_im;
  reg        [23:0]   shift_reg_863_re;
  reg        [23:0]   shift_reg_863_im;
  reg        [23:0]   shift_reg_864_re;
  reg        [23:0]   shift_reg_864_im;
  reg        [23:0]   shift_reg_865_re;
  reg        [23:0]   shift_reg_865_im;
  reg        [23:0]   shift_reg_866_re;
  reg        [23:0]   shift_reg_866_im;
  reg        [23:0]   shift_reg_867_re;
  reg        [23:0]   shift_reg_867_im;
  reg        [23:0]   shift_reg_868_re;
  reg        [23:0]   shift_reg_868_im;
  reg        [23:0]   shift_reg_869_re;
  reg        [23:0]   shift_reg_869_im;
  reg        [23:0]   shift_reg_870_re;
  reg        [23:0]   shift_reg_870_im;
  reg        [23:0]   shift_reg_871_re;
  reg        [23:0]   shift_reg_871_im;
  reg        [23:0]   shift_reg_872_re;
  reg        [23:0]   shift_reg_872_im;
  reg        [23:0]   shift_reg_873_re;
  reg        [23:0]   shift_reg_873_im;
  reg        [23:0]   shift_reg_874_re;
  reg        [23:0]   shift_reg_874_im;
  reg        [23:0]   shift_reg_875_re;
  reg        [23:0]   shift_reg_875_im;
  reg        [23:0]   shift_reg_876_re;
  reg        [23:0]   shift_reg_876_im;
  reg        [23:0]   shift_reg_877_re;
  reg        [23:0]   shift_reg_877_im;
  reg        [23:0]   shift_reg_878_re;
  reg        [23:0]   shift_reg_878_im;
  reg        [23:0]   shift_reg_879_re;
  reg        [23:0]   shift_reg_879_im;
  reg        [23:0]   shift_reg_880_re;
  reg        [23:0]   shift_reg_880_im;
  reg        [23:0]   shift_reg_881_re;
  reg        [23:0]   shift_reg_881_im;
  reg        [23:0]   shift_reg_882_re;
  reg        [23:0]   shift_reg_882_im;
  reg        [23:0]   shift_reg_883_re;
  reg        [23:0]   shift_reg_883_im;
  reg        [23:0]   shift_reg_884_re;
  reg        [23:0]   shift_reg_884_im;
  reg        [23:0]   shift_reg_885_re;
  reg        [23:0]   shift_reg_885_im;
  reg        [23:0]   shift_reg_886_re;
  reg        [23:0]   shift_reg_886_im;
  reg        [23:0]   shift_reg_887_re;
  reg        [23:0]   shift_reg_887_im;
  reg        [23:0]   shift_reg_888_re;
  reg        [23:0]   shift_reg_888_im;
  reg        [23:0]   shift_reg_889_re;
  reg        [23:0]   shift_reg_889_im;
  reg        [23:0]   shift_reg_890_re;
  reg        [23:0]   shift_reg_890_im;
  reg        [23:0]   shift_reg_891_re;
  reg        [23:0]   shift_reg_891_im;
  reg        [23:0]   shift_reg_892_re;
  reg        [23:0]   shift_reg_892_im;
  reg        [23:0]   shift_reg_893_re;
  reg        [23:0]   shift_reg_893_im;
  reg        [23:0]   shift_reg_894_re;
  reg        [23:0]   shift_reg_894_im;
  reg        [23:0]   shift_reg_895_re;
  reg        [23:0]   shift_reg_895_im;
  reg        [23:0]   shift_reg_896_re;
  reg        [23:0]   shift_reg_896_im;
  reg        [23:0]   shift_reg_897_re;
  reg        [23:0]   shift_reg_897_im;
  reg        [23:0]   shift_reg_898_re;
  reg        [23:0]   shift_reg_898_im;
  reg        [23:0]   shift_reg_899_re;
  reg        [23:0]   shift_reg_899_im;
  reg        [23:0]   shift_reg_900_re;
  reg        [23:0]   shift_reg_900_im;
  reg        [23:0]   shift_reg_901_re;
  reg        [23:0]   shift_reg_901_im;
  reg        [23:0]   shift_reg_902_re;
  reg        [23:0]   shift_reg_902_im;
  reg        [23:0]   shift_reg_903_re;
  reg        [23:0]   shift_reg_903_im;
  reg        [23:0]   shift_reg_904_re;
  reg        [23:0]   shift_reg_904_im;
  reg        [23:0]   shift_reg_905_re;
  reg        [23:0]   shift_reg_905_im;
  reg        [23:0]   shift_reg_906_re;
  reg        [23:0]   shift_reg_906_im;
  reg        [23:0]   shift_reg_907_re;
  reg        [23:0]   shift_reg_907_im;
  reg        [23:0]   shift_reg_908_re;
  reg        [23:0]   shift_reg_908_im;
  reg        [23:0]   shift_reg_909_re;
  reg        [23:0]   shift_reg_909_im;
  reg        [23:0]   shift_reg_910_re;
  reg        [23:0]   shift_reg_910_im;
  reg        [23:0]   shift_reg_911_re;
  reg        [23:0]   shift_reg_911_im;
  reg        [23:0]   shift_reg_912_re;
  reg        [23:0]   shift_reg_912_im;
  reg        [23:0]   shift_reg_913_re;
  reg        [23:0]   shift_reg_913_im;
  reg        [23:0]   shift_reg_914_re;
  reg        [23:0]   shift_reg_914_im;
  reg        [23:0]   shift_reg_915_re;
  reg        [23:0]   shift_reg_915_im;
  reg        [23:0]   shift_reg_916_re;
  reg        [23:0]   shift_reg_916_im;
  reg        [23:0]   shift_reg_917_re;
  reg        [23:0]   shift_reg_917_im;
  reg        [23:0]   shift_reg_918_re;
  reg        [23:0]   shift_reg_918_im;
  reg        [23:0]   shift_reg_919_re;
  reg        [23:0]   shift_reg_919_im;
  reg        [23:0]   shift_reg_920_re;
  reg        [23:0]   shift_reg_920_im;
  reg        [23:0]   shift_reg_921_re;
  reg        [23:0]   shift_reg_921_im;
  reg        [23:0]   shift_reg_922_re;
  reg        [23:0]   shift_reg_922_im;
  reg        [23:0]   shift_reg_923_re;
  reg        [23:0]   shift_reg_923_im;
  reg        [23:0]   shift_reg_924_re;
  reg        [23:0]   shift_reg_924_im;
  reg        [23:0]   shift_reg_925_re;
  reg        [23:0]   shift_reg_925_im;
  reg        [23:0]   shift_reg_926_re;
  reg        [23:0]   shift_reg_926_im;
  reg        [23:0]   shift_reg_927_re;
  reg        [23:0]   shift_reg_927_im;
  reg        [23:0]   shift_reg_928_re;
  reg        [23:0]   shift_reg_928_im;
  reg        [23:0]   shift_reg_929_re;
  reg        [23:0]   shift_reg_929_im;
  reg        [23:0]   shift_reg_930_re;
  reg        [23:0]   shift_reg_930_im;
  reg        [23:0]   shift_reg_931_re;
  reg        [23:0]   shift_reg_931_im;
  reg        [23:0]   shift_reg_932_re;
  reg        [23:0]   shift_reg_932_im;
  reg        [23:0]   shift_reg_933_re;
  reg        [23:0]   shift_reg_933_im;
  reg        [23:0]   shift_reg_934_re;
  reg        [23:0]   shift_reg_934_im;
  reg        [23:0]   shift_reg_935_re;
  reg        [23:0]   shift_reg_935_im;
  reg        [23:0]   shift_reg_936_re;
  reg        [23:0]   shift_reg_936_im;
  reg        [23:0]   shift_reg_937_re;
  reg        [23:0]   shift_reg_937_im;
  reg        [23:0]   shift_reg_938_re;
  reg        [23:0]   shift_reg_938_im;
  reg        [23:0]   shift_reg_939_re;
  reg        [23:0]   shift_reg_939_im;
  reg        [23:0]   shift_reg_940_re;
  reg        [23:0]   shift_reg_940_im;
  reg        [23:0]   shift_reg_941_re;
  reg        [23:0]   shift_reg_941_im;
  reg        [23:0]   shift_reg_942_re;
  reg        [23:0]   shift_reg_942_im;
  reg        [23:0]   shift_reg_943_re;
  reg        [23:0]   shift_reg_943_im;
  reg        [23:0]   shift_reg_944_re;
  reg        [23:0]   shift_reg_944_im;
  reg        [23:0]   shift_reg_945_re;
  reg        [23:0]   shift_reg_945_im;
  reg        [23:0]   shift_reg_946_re;
  reg        [23:0]   shift_reg_946_im;
  reg        [23:0]   shift_reg_947_re;
  reg        [23:0]   shift_reg_947_im;
  reg        [23:0]   shift_reg_948_re;
  reg        [23:0]   shift_reg_948_im;
  reg        [23:0]   shift_reg_949_re;
  reg        [23:0]   shift_reg_949_im;
  reg        [23:0]   shift_reg_950_re;
  reg        [23:0]   shift_reg_950_im;
  reg        [23:0]   shift_reg_951_re;
  reg        [23:0]   shift_reg_951_im;
  reg        [23:0]   shift_reg_952_re;
  reg        [23:0]   shift_reg_952_im;
  reg        [23:0]   shift_reg_953_re;
  reg        [23:0]   shift_reg_953_im;
  reg        [23:0]   shift_reg_954_re;
  reg        [23:0]   shift_reg_954_im;
  reg        [23:0]   shift_reg_955_re;
  reg        [23:0]   shift_reg_955_im;
  reg        [23:0]   shift_reg_956_re;
  reg        [23:0]   shift_reg_956_im;
  reg        [23:0]   shift_reg_957_re;
  reg        [23:0]   shift_reg_957_im;
  reg        [23:0]   shift_reg_958_re;
  reg        [23:0]   shift_reg_958_im;
  reg        [23:0]   shift_reg_959_re;
  reg        [23:0]   shift_reg_959_im;
  reg        [23:0]   shift_reg_960_re;
  reg        [23:0]   shift_reg_960_im;
  reg        [23:0]   shift_reg_961_re;
  reg        [23:0]   shift_reg_961_im;
  reg        [23:0]   shift_reg_962_re;
  reg        [23:0]   shift_reg_962_im;
  reg        [23:0]   shift_reg_963_re;
  reg        [23:0]   shift_reg_963_im;
  reg        [23:0]   shift_reg_964_re;
  reg        [23:0]   shift_reg_964_im;
  reg        [23:0]   shift_reg_965_re;
  reg        [23:0]   shift_reg_965_im;
  reg        [23:0]   shift_reg_966_re;
  reg        [23:0]   shift_reg_966_im;
  reg        [23:0]   shift_reg_967_re;
  reg        [23:0]   shift_reg_967_im;
  reg        [23:0]   shift_reg_968_re;
  reg        [23:0]   shift_reg_968_im;
  reg        [23:0]   shift_reg_969_re;
  reg        [23:0]   shift_reg_969_im;
  reg        [23:0]   shift_reg_970_re;
  reg        [23:0]   shift_reg_970_im;
  reg        [23:0]   shift_reg_971_re;
  reg        [23:0]   shift_reg_971_im;
  reg        [23:0]   shift_reg_972_re;
  reg        [23:0]   shift_reg_972_im;
  reg        [23:0]   shift_reg_973_re;
  reg        [23:0]   shift_reg_973_im;
  reg        [23:0]   shift_reg_974_re;
  reg        [23:0]   shift_reg_974_im;
  reg        [23:0]   shift_reg_975_re;
  reg        [23:0]   shift_reg_975_im;
  reg        [23:0]   shift_reg_976_re;
  reg        [23:0]   shift_reg_976_im;
  reg        [23:0]   shift_reg_977_re;
  reg        [23:0]   shift_reg_977_im;
  reg        [23:0]   shift_reg_978_re;
  reg        [23:0]   shift_reg_978_im;
  reg        [23:0]   shift_reg_979_re;
  reg        [23:0]   shift_reg_979_im;
  reg        [23:0]   shift_reg_980_re;
  reg        [23:0]   shift_reg_980_im;
  reg        [23:0]   shift_reg_981_re;
  reg        [23:0]   shift_reg_981_im;
  reg        [23:0]   shift_reg_982_re;
  reg        [23:0]   shift_reg_982_im;
  reg        [23:0]   shift_reg_983_re;
  reg        [23:0]   shift_reg_983_im;
  reg        [23:0]   shift_reg_984_re;
  reg        [23:0]   shift_reg_984_im;
  reg        [23:0]   shift_reg_985_re;
  reg        [23:0]   shift_reg_985_im;
  reg        [23:0]   shift_reg_986_re;
  reg        [23:0]   shift_reg_986_im;
  reg        [23:0]   shift_reg_987_re;
  reg        [23:0]   shift_reg_987_im;
  reg        [23:0]   shift_reg_988_re;
  reg        [23:0]   shift_reg_988_im;
  reg        [23:0]   shift_reg_989_re;
  reg        [23:0]   shift_reg_989_im;
  reg        [23:0]   shift_reg_990_re;
  reg        [23:0]   shift_reg_990_im;
  reg        [23:0]   shift_reg_991_re;
  reg        [23:0]   shift_reg_991_im;
  reg        [23:0]   shift_reg_992_re;
  reg        [23:0]   shift_reg_992_im;
  reg        [23:0]   shift_reg_993_re;
  reg        [23:0]   shift_reg_993_im;
  reg        [23:0]   shift_reg_994_re;
  reg        [23:0]   shift_reg_994_im;
  reg        [23:0]   shift_reg_995_re;
  reg        [23:0]   shift_reg_995_im;
  reg        [23:0]   shift_reg_996_re;
  reg        [23:0]   shift_reg_996_im;
  reg        [23:0]   shift_reg_997_re;
  reg        [23:0]   shift_reg_997_im;
  reg        [23:0]   shift_reg_998_re;
  reg        [23:0]   shift_reg_998_im;
  reg        [23:0]   shift_reg_999_re;
  reg        [23:0]   shift_reg_999_im;
  reg        [23:0]   shift_reg_1000_re;
  reg        [23:0]   shift_reg_1000_im;
  reg        [23:0]   shift_reg_1001_re;
  reg        [23:0]   shift_reg_1001_im;
  reg        [23:0]   shift_reg_1002_re;
  reg        [23:0]   shift_reg_1002_im;
  reg        [23:0]   shift_reg_1003_re;
  reg        [23:0]   shift_reg_1003_im;
  reg        [23:0]   shift_reg_1004_re;
  reg        [23:0]   shift_reg_1004_im;
  reg        [23:0]   shift_reg_1005_re;
  reg        [23:0]   shift_reg_1005_im;
  reg        [23:0]   shift_reg_1006_re;
  reg        [23:0]   shift_reg_1006_im;
  reg        [23:0]   shift_reg_1007_re;
  reg        [23:0]   shift_reg_1007_im;
  reg        [23:0]   shift_reg_1008_re;
  reg        [23:0]   shift_reg_1008_im;
  reg        [23:0]   shift_reg_1009_re;
  reg        [23:0]   shift_reg_1009_im;
  reg        [23:0]   shift_reg_1010_re;
  reg        [23:0]   shift_reg_1010_im;
  reg        [23:0]   shift_reg_1011_re;
  reg        [23:0]   shift_reg_1011_im;
  reg        [23:0]   shift_reg_1012_re;
  reg        [23:0]   shift_reg_1012_im;
  reg        [23:0]   shift_reg_1013_re;
  reg        [23:0]   shift_reg_1013_im;
  reg        [23:0]   shift_reg_1014_re;
  reg        [23:0]   shift_reg_1014_im;
  reg        [23:0]   shift_reg_1015_re;
  reg        [23:0]   shift_reg_1015_im;
  reg        [23:0]   shift_reg_1016_re;
  reg        [23:0]   shift_reg_1016_im;
  reg        [23:0]   shift_reg_1017_re;
  reg        [23:0]   shift_reg_1017_im;
  reg        [23:0]   shift_reg_1018_re;
  reg        [23:0]   shift_reg_1018_im;
  reg        [23:0]   shift_reg_1019_re;
  reg        [23:0]   shift_reg_1019_im;
  reg        [23:0]   shift_reg_1020_re;
  reg        [23:0]   shift_reg_1020_im;
  reg        [23:0]   shift_reg_1021_re;
  reg        [23:0]   shift_reg_1021_im;
  reg        [23:0]   shift_reg_1022_re;
  reg        [23:0]   shift_reg_1022_im;
  reg        [23:0]   shift_reg_1023_re;
  reg        [23:0]   shift_reg_1023_im;

  assign output_re = shift_reg_1023_re;
  assign output_im = shift_reg_1023_im;
  always @(posedge clk) begin
    shift_reg_0_re <= input_re;
    shift_reg_0_im <= input_im;
    shift_reg_1_re <= shift_reg_0_re;
    shift_reg_1_im <= shift_reg_0_im;
    shift_reg_2_re <= shift_reg_1_re;
    shift_reg_2_im <= shift_reg_1_im;
    shift_reg_3_re <= shift_reg_2_re;
    shift_reg_3_im <= shift_reg_2_im;
    shift_reg_4_re <= shift_reg_3_re;
    shift_reg_4_im <= shift_reg_3_im;
    shift_reg_5_re <= shift_reg_4_re;
    shift_reg_5_im <= shift_reg_4_im;
    shift_reg_6_re <= shift_reg_5_re;
    shift_reg_6_im <= shift_reg_5_im;
    shift_reg_7_re <= shift_reg_6_re;
    shift_reg_7_im <= shift_reg_6_im;
    shift_reg_8_re <= shift_reg_7_re;
    shift_reg_8_im <= shift_reg_7_im;
    shift_reg_9_re <= shift_reg_8_re;
    shift_reg_9_im <= shift_reg_8_im;
    shift_reg_10_re <= shift_reg_9_re;
    shift_reg_10_im <= shift_reg_9_im;
    shift_reg_11_re <= shift_reg_10_re;
    shift_reg_11_im <= shift_reg_10_im;
    shift_reg_12_re <= shift_reg_11_re;
    shift_reg_12_im <= shift_reg_11_im;
    shift_reg_13_re <= shift_reg_12_re;
    shift_reg_13_im <= shift_reg_12_im;
    shift_reg_14_re <= shift_reg_13_re;
    shift_reg_14_im <= shift_reg_13_im;
    shift_reg_15_re <= shift_reg_14_re;
    shift_reg_15_im <= shift_reg_14_im;
    shift_reg_16_re <= shift_reg_15_re;
    shift_reg_16_im <= shift_reg_15_im;
    shift_reg_17_re <= shift_reg_16_re;
    shift_reg_17_im <= shift_reg_16_im;
    shift_reg_18_re <= shift_reg_17_re;
    shift_reg_18_im <= shift_reg_17_im;
    shift_reg_19_re <= shift_reg_18_re;
    shift_reg_19_im <= shift_reg_18_im;
    shift_reg_20_re <= shift_reg_19_re;
    shift_reg_20_im <= shift_reg_19_im;
    shift_reg_21_re <= shift_reg_20_re;
    shift_reg_21_im <= shift_reg_20_im;
    shift_reg_22_re <= shift_reg_21_re;
    shift_reg_22_im <= shift_reg_21_im;
    shift_reg_23_re <= shift_reg_22_re;
    shift_reg_23_im <= shift_reg_22_im;
    shift_reg_24_re <= shift_reg_23_re;
    shift_reg_24_im <= shift_reg_23_im;
    shift_reg_25_re <= shift_reg_24_re;
    shift_reg_25_im <= shift_reg_24_im;
    shift_reg_26_re <= shift_reg_25_re;
    shift_reg_26_im <= shift_reg_25_im;
    shift_reg_27_re <= shift_reg_26_re;
    shift_reg_27_im <= shift_reg_26_im;
    shift_reg_28_re <= shift_reg_27_re;
    shift_reg_28_im <= shift_reg_27_im;
    shift_reg_29_re <= shift_reg_28_re;
    shift_reg_29_im <= shift_reg_28_im;
    shift_reg_30_re <= shift_reg_29_re;
    shift_reg_30_im <= shift_reg_29_im;
    shift_reg_31_re <= shift_reg_30_re;
    shift_reg_31_im <= shift_reg_30_im;
    shift_reg_32_re <= shift_reg_31_re;
    shift_reg_32_im <= shift_reg_31_im;
    shift_reg_33_re <= shift_reg_32_re;
    shift_reg_33_im <= shift_reg_32_im;
    shift_reg_34_re <= shift_reg_33_re;
    shift_reg_34_im <= shift_reg_33_im;
    shift_reg_35_re <= shift_reg_34_re;
    shift_reg_35_im <= shift_reg_34_im;
    shift_reg_36_re <= shift_reg_35_re;
    shift_reg_36_im <= shift_reg_35_im;
    shift_reg_37_re <= shift_reg_36_re;
    shift_reg_37_im <= shift_reg_36_im;
    shift_reg_38_re <= shift_reg_37_re;
    shift_reg_38_im <= shift_reg_37_im;
    shift_reg_39_re <= shift_reg_38_re;
    shift_reg_39_im <= shift_reg_38_im;
    shift_reg_40_re <= shift_reg_39_re;
    shift_reg_40_im <= shift_reg_39_im;
    shift_reg_41_re <= shift_reg_40_re;
    shift_reg_41_im <= shift_reg_40_im;
    shift_reg_42_re <= shift_reg_41_re;
    shift_reg_42_im <= shift_reg_41_im;
    shift_reg_43_re <= shift_reg_42_re;
    shift_reg_43_im <= shift_reg_42_im;
    shift_reg_44_re <= shift_reg_43_re;
    shift_reg_44_im <= shift_reg_43_im;
    shift_reg_45_re <= shift_reg_44_re;
    shift_reg_45_im <= shift_reg_44_im;
    shift_reg_46_re <= shift_reg_45_re;
    shift_reg_46_im <= shift_reg_45_im;
    shift_reg_47_re <= shift_reg_46_re;
    shift_reg_47_im <= shift_reg_46_im;
    shift_reg_48_re <= shift_reg_47_re;
    shift_reg_48_im <= shift_reg_47_im;
    shift_reg_49_re <= shift_reg_48_re;
    shift_reg_49_im <= shift_reg_48_im;
    shift_reg_50_re <= shift_reg_49_re;
    shift_reg_50_im <= shift_reg_49_im;
    shift_reg_51_re <= shift_reg_50_re;
    shift_reg_51_im <= shift_reg_50_im;
    shift_reg_52_re <= shift_reg_51_re;
    shift_reg_52_im <= shift_reg_51_im;
    shift_reg_53_re <= shift_reg_52_re;
    shift_reg_53_im <= shift_reg_52_im;
    shift_reg_54_re <= shift_reg_53_re;
    shift_reg_54_im <= shift_reg_53_im;
    shift_reg_55_re <= shift_reg_54_re;
    shift_reg_55_im <= shift_reg_54_im;
    shift_reg_56_re <= shift_reg_55_re;
    shift_reg_56_im <= shift_reg_55_im;
    shift_reg_57_re <= shift_reg_56_re;
    shift_reg_57_im <= shift_reg_56_im;
    shift_reg_58_re <= shift_reg_57_re;
    shift_reg_58_im <= shift_reg_57_im;
    shift_reg_59_re <= shift_reg_58_re;
    shift_reg_59_im <= shift_reg_58_im;
    shift_reg_60_re <= shift_reg_59_re;
    shift_reg_60_im <= shift_reg_59_im;
    shift_reg_61_re <= shift_reg_60_re;
    shift_reg_61_im <= shift_reg_60_im;
    shift_reg_62_re <= shift_reg_61_re;
    shift_reg_62_im <= shift_reg_61_im;
    shift_reg_63_re <= shift_reg_62_re;
    shift_reg_63_im <= shift_reg_62_im;
    shift_reg_64_re <= shift_reg_63_re;
    shift_reg_64_im <= shift_reg_63_im;
    shift_reg_65_re <= shift_reg_64_re;
    shift_reg_65_im <= shift_reg_64_im;
    shift_reg_66_re <= shift_reg_65_re;
    shift_reg_66_im <= shift_reg_65_im;
    shift_reg_67_re <= shift_reg_66_re;
    shift_reg_67_im <= shift_reg_66_im;
    shift_reg_68_re <= shift_reg_67_re;
    shift_reg_68_im <= shift_reg_67_im;
    shift_reg_69_re <= shift_reg_68_re;
    shift_reg_69_im <= shift_reg_68_im;
    shift_reg_70_re <= shift_reg_69_re;
    shift_reg_70_im <= shift_reg_69_im;
    shift_reg_71_re <= shift_reg_70_re;
    shift_reg_71_im <= shift_reg_70_im;
    shift_reg_72_re <= shift_reg_71_re;
    shift_reg_72_im <= shift_reg_71_im;
    shift_reg_73_re <= shift_reg_72_re;
    shift_reg_73_im <= shift_reg_72_im;
    shift_reg_74_re <= shift_reg_73_re;
    shift_reg_74_im <= shift_reg_73_im;
    shift_reg_75_re <= shift_reg_74_re;
    shift_reg_75_im <= shift_reg_74_im;
    shift_reg_76_re <= shift_reg_75_re;
    shift_reg_76_im <= shift_reg_75_im;
    shift_reg_77_re <= shift_reg_76_re;
    shift_reg_77_im <= shift_reg_76_im;
    shift_reg_78_re <= shift_reg_77_re;
    shift_reg_78_im <= shift_reg_77_im;
    shift_reg_79_re <= shift_reg_78_re;
    shift_reg_79_im <= shift_reg_78_im;
    shift_reg_80_re <= shift_reg_79_re;
    shift_reg_80_im <= shift_reg_79_im;
    shift_reg_81_re <= shift_reg_80_re;
    shift_reg_81_im <= shift_reg_80_im;
    shift_reg_82_re <= shift_reg_81_re;
    shift_reg_82_im <= shift_reg_81_im;
    shift_reg_83_re <= shift_reg_82_re;
    shift_reg_83_im <= shift_reg_82_im;
    shift_reg_84_re <= shift_reg_83_re;
    shift_reg_84_im <= shift_reg_83_im;
    shift_reg_85_re <= shift_reg_84_re;
    shift_reg_85_im <= shift_reg_84_im;
    shift_reg_86_re <= shift_reg_85_re;
    shift_reg_86_im <= shift_reg_85_im;
    shift_reg_87_re <= shift_reg_86_re;
    shift_reg_87_im <= shift_reg_86_im;
    shift_reg_88_re <= shift_reg_87_re;
    shift_reg_88_im <= shift_reg_87_im;
    shift_reg_89_re <= shift_reg_88_re;
    shift_reg_89_im <= shift_reg_88_im;
    shift_reg_90_re <= shift_reg_89_re;
    shift_reg_90_im <= shift_reg_89_im;
    shift_reg_91_re <= shift_reg_90_re;
    shift_reg_91_im <= shift_reg_90_im;
    shift_reg_92_re <= shift_reg_91_re;
    shift_reg_92_im <= shift_reg_91_im;
    shift_reg_93_re <= shift_reg_92_re;
    shift_reg_93_im <= shift_reg_92_im;
    shift_reg_94_re <= shift_reg_93_re;
    shift_reg_94_im <= shift_reg_93_im;
    shift_reg_95_re <= shift_reg_94_re;
    shift_reg_95_im <= shift_reg_94_im;
    shift_reg_96_re <= shift_reg_95_re;
    shift_reg_96_im <= shift_reg_95_im;
    shift_reg_97_re <= shift_reg_96_re;
    shift_reg_97_im <= shift_reg_96_im;
    shift_reg_98_re <= shift_reg_97_re;
    shift_reg_98_im <= shift_reg_97_im;
    shift_reg_99_re <= shift_reg_98_re;
    shift_reg_99_im <= shift_reg_98_im;
    shift_reg_100_re <= shift_reg_99_re;
    shift_reg_100_im <= shift_reg_99_im;
    shift_reg_101_re <= shift_reg_100_re;
    shift_reg_101_im <= shift_reg_100_im;
    shift_reg_102_re <= shift_reg_101_re;
    shift_reg_102_im <= shift_reg_101_im;
    shift_reg_103_re <= shift_reg_102_re;
    shift_reg_103_im <= shift_reg_102_im;
    shift_reg_104_re <= shift_reg_103_re;
    shift_reg_104_im <= shift_reg_103_im;
    shift_reg_105_re <= shift_reg_104_re;
    shift_reg_105_im <= shift_reg_104_im;
    shift_reg_106_re <= shift_reg_105_re;
    shift_reg_106_im <= shift_reg_105_im;
    shift_reg_107_re <= shift_reg_106_re;
    shift_reg_107_im <= shift_reg_106_im;
    shift_reg_108_re <= shift_reg_107_re;
    shift_reg_108_im <= shift_reg_107_im;
    shift_reg_109_re <= shift_reg_108_re;
    shift_reg_109_im <= shift_reg_108_im;
    shift_reg_110_re <= shift_reg_109_re;
    shift_reg_110_im <= shift_reg_109_im;
    shift_reg_111_re <= shift_reg_110_re;
    shift_reg_111_im <= shift_reg_110_im;
    shift_reg_112_re <= shift_reg_111_re;
    shift_reg_112_im <= shift_reg_111_im;
    shift_reg_113_re <= shift_reg_112_re;
    shift_reg_113_im <= shift_reg_112_im;
    shift_reg_114_re <= shift_reg_113_re;
    shift_reg_114_im <= shift_reg_113_im;
    shift_reg_115_re <= shift_reg_114_re;
    shift_reg_115_im <= shift_reg_114_im;
    shift_reg_116_re <= shift_reg_115_re;
    shift_reg_116_im <= shift_reg_115_im;
    shift_reg_117_re <= shift_reg_116_re;
    shift_reg_117_im <= shift_reg_116_im;
    shift_reg_118_re <= shift_reg_117_re;
    shift_reg_118_im <= shift_reg_117_im;
    shift_reg_119_re <= shift_reg_118_re;
    shift_reg_119_im <= shift_reg_118_im;
    shift_reg_120_re <= shift_reg_119_re;
    shift_reg_120_im <= shift_reg_119_im;
    shift_reg_121_re <= shift_reg_120_re;
    shift_reg_121_im <= shift_reg_120_im;
    shift_reg_122_re <= shift_reg_121_re;
    shift_reg_122_im <= shift_reg_121_im;
    shift_reg_123_re <= shift_reg_122_re;
    shift_reg_123_im <= shift_reg_122_im;
    shift_reg_124_re <= shift_reg_123_re;
    shift_reg_124_im <= shift_reg_123_im;
    shift_reg_125_re <= shift_reg_124_re;
    shift_reg_125_im <= shift_reg_124_im;
    shift_reg_126_re <= shift_reg_125_re;
    shift_reg_126_im <= shift_reg_125_im;
    shift_reg_127_re <= shift_reg_126_re;
    shift_reg_127_im <= shift_reg_126_im;
    shift_reg_128_re <= shift_reg_127_re;
    shift_reg_128_im <= shift_reg_127_im;
    shift_reg_129_re <= shift_reg_128_re;
    shift_reg_129_im <= shift_reg_128_im;
    shift_reg_130_re <= shift_reg_129_re;
    shift_reg_130_im <= shift_reg_129_im;
    shift_reg_131_re <= shift_reg_130_re;
    shift_reg_131_im <= shift_reg_130_im;
    shift_reg_132_re <= shift_reg_131_re;
    shift_reg_132_im <= shift_reg_131_im;
    shift_reg_133_re <= shift_reg_132_re;
    shift_reg_133_im <= shift_reg_132_im;
    shift_reg_134_re <= shift_reg_133_re;
    shift_reg_134_im <= shift_reg_133_im;
    shift_reg_135_re <= shift_reg_134_re;
    shift_reg_135_im <= shift_reg_134_im;
    shift_reg_136_re <= shift_reg_135_re;
    shift_reg_136_im <= shift_reg_135_im;
    shift_reg_137_re <= shift_reg_136_re;
    shift_reg_137_im <= shift_reg_136_im;
    shift_reg_138_re <= shift_reg_137_re;
    shift_reg_138_im <= shift_reg_137_im;
    shift_reg_139_re <= shift_reg_138_re;
    shift_reg_139_im <= shift_reg_138_im;
    shift_reg_140_re <= shift_reg_139_re;
    shift_reg_140_im <= shift_reg_139_im;
    shift_reg_141_re <= shift_reg_140_re;
    shift_reg_141_im <= shift_reg_140_im;
    shift_reg_142_re <= shift_reg_141_re;
    shift_reg_142_im <= shift_reg_141_im;
    shift_reg_143_re <= shift_reg_142_re;
    shift_reg_143_im <= shift_reg_142_im;
    shift_reg_144_re <= shift_reg_143_re;
    shift_reg_144_im <= shift_reg_143_im;
    shift_reg_145_re <= shift_reg_144_re;
    shift_reg_145_im <= shift_reg_144_im;
    shift_reg_146_re <= shift_reg_145_re;
    shift_reg_146_im <= shift_reg_145_im;
    shift_reg_147_re <= shift_reg_146_re;
    shift_reg_147_im <= shift_reg_146_im;
    shift_reg_148_re <= shift_reg_147_re;
    shift_reg_148_im <= shift_reg_147_im;
    shift_reg_149_re <= shift_reg_148_re;
    shift_reg_149_im <= shift_reg_148_im;
    shift_reg_150_re <= shift_reg_149_re;
    shift_reg_150_im <= shift_reg_149_im;
    shift_reg_151_re <= shift_reg_150_re;
    shift_reg_151_im <= shift_reg_150_im;
    shift_reg_152_re <= shift_reg_151_re;
    shift_reg_152_im <= shift_reg_151_im;
    shift_reg_153_re <= shift_reg_152_re;
    shift_reg_153_im <= shift_reg_152_im;
    shift_reg_154_re <= shift_reg_153_re;
    shift_reg_154_im <= shift_reg_153_im;
    shift_reg_155_re <= shift_reg_154_re;
    shift_reg_155_im <= shift_reg_154_im;
    shift_reg_156_re <= shift_reg_155_re;
    shift_reg_156_im <= shift_reg_155_im;
    shift_reg_157_re <= shift_reg_156_re;
    shift_reg_157_im <= shift_reg_156_im;
    shift_reg_158_re <= shift_reg_157_re;
    shift_reg_158_im <= shift_reg_157_im;
    shift_reg_159_re <= shift_reg_158_re;
    shift_reg_159_im <= shift_reg_158_im;
    shift_reg_160_re <= shift_reg_159_re;
    shift_reg_160_im <= shift_reg_159_im;
    shift_reg_161_re <= shift_reg_160_re;
    shift_reg_161_im <= shift_reg_160_im;
    shift_reg_162_re <= shift_reg_161_re;
    shift_reg_162_im <= shift_reg_161_im;
    shift_reg_163_re <= shift_reg_162_re;
    shift_reg_163_im <= shift_reg_162_im;
    shift_reg_164_re <= shift_reg_163_re;
    shift_reg_164_im <= shift_reg_163_im;
    shift_reg_165_re <= shift_reg_164_re;
    shift_reg_165_im <= shift_reg_164_im;
    shift_reg_166_re <= shift_reg_165_re;
    shift_reg_166_im <= shift_reg_165_im;
    shift_reg_167_re <= shift_reg_166_re;
    shift_reg_167_im <= shift_reg_166_im;
    shift_reg_168_re <= shift_reg_167_re;
    shift_reg_168_im <= shift_reg_167_im;
    shift_reg_169_re <= shift_reg_168_re;
    shift_reg_169_im <= shift_reg_168_im;
    shift_reg_170_re <= shift_reg_169_re;
    shift_reg_170_im <= shift_reg_169_im;
    shift_reg_171_re <= shift_reg_170_re;
    shift_reg_171_im <= shift_reg_170_im;
    shift_reg_172_re <= shift_reg_171_re;
    shift_reg_172_im <= shift_reg_171_im;
    shift_reg_173_re <= shift_reg_172_re;
    shift_reg_173_im <= shift_reg_172_im;
    shift_reg_174_re <= shift_reg_173_re;
    shift_reg_174_im <= shift_reg_173_im;
    shift_reg_175_re <= shift_reg_174_re;
    shift_reg_175_im <= shift_reg_174_im;
    shift_reg_176_re <= shift_reg_175_re;
    shift_reg_176_im <= shift_reg_175_im;
    shift_reg_177_re <= shift_reg_176_re;
    shift_reg_177_im <= shift_reg_176_im;
    shift_reg_178_re <= shift_reg_177_re;
    shift_reg_178_im <= shift_reg_177_im;
    shift_reg_179_re <= shift_reg_178_re;
    shift_reg_179_im <= shift_reg_178_im;
    shift_reg_180_re <= shift_reg_179_re;
    shift_reg_180_im <= shift_reg_179_im;
    shift_reg_181_re <= shift_reg_180_re;
    shift_reg_181_im <= shift_reg_180_im;
    shift_reg_182_re <= shift_reg_181_re;
    shift_reg_182_im <= shift_reg_181_im;
    shift_reg_183_re <= shift_reg_182_re;
    shift_reg_183_im <= shift_reg_182_im;
    shift_reg_184_re <= shift_reg_183_re;
    shift_reg_184_im <= shift_reg_183_im;
    shift_reg_185_re <= shift_reg_184_re;
    shift_reg_185_im <= shift_reg_184_im;
    shift_reg_186_re <= shift_reg_185_re;
    shift_reg_186_im <= shift_reg_185_im;
    shift_reg_187_re <= shift_reg_186_re;
    shift_reg_187_im <= shift_reg_186_im;
    shift_reg_188_re <= shift_reg_187_re;
    shift_reg_188_im <= shift_reg_187_im;
    shift_reg_189_re <= shift_reg_188_re;
    shift_reg_189_im <= shift_reg_188_im;
    shift_reg_190_re <= shift_reg_189_re;
    shift_reg_190_im <= shift_reg_189_im;
    shift_reg_191_re <= shift_reg_190_re;
    shift_reg_191_im <= shift_reg_190_im;
    shift_reg_192_re <= shift_reg_191_re;
    shift_reg_192_im <= shift_reg_191_im;
    shift_reg_193_re <= shift_reg_192_re;
    shift_reg_193_im <= shift_reg_192_im;
    shift_reg_194_re <= shift_reg_193_re;
    shift_reg_194_im <= shift_reg_193_im;
    shift_reg_195_re <= shift_reg_194_re;
    shift_reg_195_im <= shift_reg_194_im;
    shift_reg_196_re <= shift_reg_195_re;
    shift_reg_196_im <= shift_reg_195_im;
    shift_reg_197_re <= shift_reg_196_re;
    shift_reg_197_im <= shift_reg_196_im;
    shift_reg_198_re <= shift_reg_197_re;
    shift_reg_198_im <= shift_reg_197_im;
    shift_reg_199_re <= shift_reg_198_re;
    shift_reg_199_im <= shift_reg_198_im;
    shift_reg_200_re <= shift_reg_199_re;
    shift_reg_200_im <= shift_reg_199_im;
    shift_reg_201_re <= shift_reg_200_re;
    shift_reg_201_im <= shift_reg_200_im;
    shift_reg_202_re <= shift_reg_201_re;
    shift_reg_202_im <= shift_reg_201_im;
    shift_reg_203_re <= shift_reg_202_re;
    shift_reg_203_im <= shift_reg_202_im;
    shift_reg_204_re <= shift_reg_203_re;
    shift_reg_204_im <= shift_reg_203_im;
    shift_reg_205_re <= shift_reg_204_re;
    shift_reg_205_im <= shift_reg_204_im;
    shift_reg_206_re <= shift_reg_205_re;
    shift_reg_206_im <= shift_reg_205_im;
    shift_reg_207_re <= shift_reg_206_re;
    shift_reg_207_im <= shift_reg_206_im;
    shift_reg_208_re <= shift_reg_207_re;
    shift_reg_208_im <= shift_reg_207_im;
    shift_reg_209_re <= shift_reg_208_re;
    shift_reg_209_im <= shift_reg_208_im;
    shift_reg_210_re <= shift_reg_209_re;
    shift_reg_210_im <= shift_reg_209_im;
    shift_reg_211_re <= shift_reg_210_re;
    shift_reg_211_im <= shift_reg_210_im;
    shift_reg_212_re <= shift_reg_211_re;
    shift_reg_212_im <= shift_reg_211_im;
    shift_reg_213_re <= shift_reg_212_re;
    shift_reg_213_im <= shift_reg_212_im;
    shift_reg_214_re <= shift_reg_213_re;
    shift_reg_214_im <= shift_reg_213_im;
    shift_reg_215_re <= shift_reg_214_re;
    shift_reg_215_im <= shift_reg_214_im;
    shift_reg_216_re <= shift_reg_215_re;
    shift_reg_216_im <= shift_reg_215_im;
    shift_reg_217_re <= shift_reg_216_re;
    shift_reg_217_im <= shift_reg_216_im;
    shift_reg_218_re <= shift_reg_217_re;
    shift_reg_218_im <= shift_reg_217_im;
    shift_reg_219_re <= shift_reg_218_re;
    shift_reg_219_im <= shift_reg_218_im;
    shift_reg_220_re <= shift_reg_219_re;
    shift_reg_220_im <= shift_reg_219_im;
    shift_reg_221_re <= shift_reg_220_re;
    shift_reg_221_im <= shift_reg_220_im;
    shift_reg_222_re <= shift_reg_221_re;
    shift_reg_222_im <= shift_reg_221_im;
    shift_reg_223_re <= shift_reg_222_re;
    shift_reg_223_im <= shift_reg_222_im;
    shift_reg_224_re <= shift_reg_223_re;
    shift_reg_224_im <= shift_reg_223_im;
    shift_reg_225_re <= shift_reg_224_re;
    shift_reg_225_im <= shift_reg_224_im;
    shift_reg_226_re <= shift_reg_225_re;
    shift_reg_226_im <= shift_reg_225_im;
    shift_reg_227_re <= shift_reg_226_re;
    shift_reg_227_im <= shift_reg_226_im;
    shift_reg_228_re <= shift_reg_227_re;
    shift_reg_228_im <= shift_reg_227_im;
    shift_reg_229_re <= shift_reg_228_re;
    shift_reg_229_im <= shift_reg_228_im;
    shift_reg_230_re <= shift_reg_229_re;
    shift_reg_230_im <= shift_reg_229_im;
    shift_reg_231_re <= shift_reg_230_re;
    shift_reg_231_im <= shift_reg_230_im;
    shift_reg_232_re <= shift_reg_231_re;
    shift_reg_232_im <= shift_reg_231_im;
    shift_reg_233_re <= shift_reg_232_re;
    shift_reg_233_im <= shift_reg_232_im;
    shift_reg_234_re <= shift_reg_233_re;
    shift_reg_234_im <= shift_reg_233_im;
    shift_reg_235_re <= shift_reg_234_re;
    shift_reg_235_im <= shift_reg_234_im;
    shift_reg_236_re <= shift_reg_235_re;
    shift_reg_236_im <= shift_reg_235_im;
    shift_reg_237_re <= shift_reg_236_re;
    shift_reg_237_im <= shift_reg_236_im;
    shift_reg_238_re <= shift_reg_237_re;
    shift_reg_238_im <= shift_reg_237_im;
    shift_reg_239_re <= shift_reg_238_re;
    shift_reg_239_im <= shift_reg_238_im;
    shift_reg_240_re <= shift_reg_239_re;
    shift_reg_240_im <= shift_reg_239_im;
    shift_reg_241_re <= shift_reg_240_re;
    shift_reg_241_im <= shift_reg_240_im;
    shift_reg_242_re <= shift_reg_241_re;
    shift_reg_242_im <= shift_reg_241_im;
    shift_reg_243_re <= shift_reg_242_re;
    shift_reg_243_im <= shift_reg_242_im;
    shift_reg_244_re <= shift_reg_243_re;
    shift_reg_244_im <= shift_reg_243_im;
    shift_reg_245_re <= shift_reg_244_re;
    shift_reg_245_im <= shift_reg_244_im;
    shift_reg_246_re <= shift_reg_245_re;
    shift_reg_246_im <= shift_reg_245_im;
    shift_reg_247_re <= shift_reg_246_re;
    shift_reg_247_im <= shift_reg_246_im;
    shift_reg_248_re <= shift_reg_247_re;
    shift_reg_248_im <= shift_reg_247_im;
    shift_reg_249_re <= shift_reg_248_re;
    shift_reg_249_im <= shift_reg_248_im;
    shift_reg_250_re <= shift_reg_249_re;
    shift_reg_250_im <= shift_reg_249_im;
    shift_reg_251_re <= shift_reg_250_re;
    shift_reg_251_im <= shift_reg_250_im;
    shift_reg_252_re <= shift_reg_251_re;
    shift_reg_252_im <= shift_reg_251_im;
    shift_reg_253_re <= shift_reg_252_re;
    shift_reg_253_im <= shift_reg_252_im;
    shift_reg_254_re <= shift_reg_253_re;
    shift_reg_254_im <= shift_reg_253_im;
    shift_reg_255_re <= shift_reg_254_re;
    shift_reg_255_im <= shift_reg_254_im;
    shift_reg_256_re <= shift_reg_255_re;
    shift_reg_256_im <= shift_reg_255_im;
    shift_reg_257_re <= shift_reg_256_re;
    shift_reg_257_im <= shift_reg_256_im;
    shift_reg_258_re <= shift_reg_257_re;
    shift_reg_258_im <= shift_reg_257_im;
    shift_reg_259_re <= shift_reg_258_re;
    shift_reg_259_im <= shift_reg_258_im;
    shift_reg_260_re <= shift_reg_259_re;
    shift_reg_260_im <= shift_reg_259_im;
    shift_reg_261_re <= shift_reg_260_re;
    shift_reg_261_im <= shift_reg_260_im;
    shift_reg_262_re <= shift_reg_261_re;
    shift_reg_262_im <= shift_reg_261_im;
    shift_reg_263_re <= shift_reg_262_re;
    shift_reg_263_im <= shift_reg_262_im;
    shift_reg_264_re <= shift_reg_263_re;
    shift_reg_264_im <= shift_reg_263_im;
    shift_reg_265_re <= shift_reg_264_re;
    shift_reg_265_im <= shift_reg_264_im;
    shift_reg_266_re <= shift_reg_265_re;
    shift_reg_266_im <= shift_reg_265_im;
    shift_reg_267_re <= shift_reg_266_re;
    shift_reg_267_im <= shift_reg_266_im;
    shift_reg_268_re <= shift_reg_267_re;
    shift_reg_268_im <= shift_reg_267_im;
    shift_reg_269_re <= shift_reg_268_re;
    shift_reg_269_im <= shift_reg_268_im;
    shift_reg_270_re <= shift_reg_269_re;
    shift_reg_270_im <= shift_reg_269_im;
    shift_reg_271_re <= shift_reg_270_re;
    shift_reg_271_im <= shift_reg_270_im;
    shift_reg_272_re <= shift_reg_271_re;
    shift_reg_272_im <= shift_reg_271_im;
    shift_reg_273_re <= shift_reg_272_re;
    shift_reg_273_im <= shift_reg_272_im;
    shift_reg_274_re <= shift_reg_273_re;
    shift_reg_274_im <= shift_reg_273_im;
    shift_reg_275_re <= shift_reg_274_re;
    shift_reg_275_im <= shift_reg_274_im;
    shift_reg_276_re <= shift_reg_275_re;
    shift_reg_276_im <= shift_reg_275_im;
    shift_reg_277_re <= shift_reg_276_re;
    shift_reg_277_im <= shift_reg_276_im;
    shift_reg_278_re <= shift_reg_277_re;
    shift_reg_278_im <= shift_reg_277_im;
    shift_reg_279_re <= shift_reg_278_re;
    shift_reg_279_im <= shift_reg_278_im;
    shift_reg_280_re <= shift_reg_279_re;
    shift_reg_280_im <= shift_reg_279_im;
    shift_reg_281_re <= shift_reg_280_re;
    shift_reg_281_im <= shift_reg_280_im;
    shift_reg_282_re <= shift_reg_281_re;
    shift_reg_282_im <= shift_reg_281_im;
    shift_reg_283_re <= shift_reg_282_re;
    shift_reg_283_im <= shift_reg_282_im;
    shift_reg_284_re <= shift_reg_283_re;
    shift_reg_284_im <= shift_reg_283_im;
    shift_reg_285_re <= shift_reg_284_re;
    shift_reg_285_im <= shift_reg_284_im;
    shift_reg_286_re <= shift_reg_285_re;
    shift_reg_286_im <= shift_reg_285_im;
    shift_reg_287_re <= shift_reg_286_re;
    shift_reg_287_im <= shift_reg_286_im;
    shift_reg_288_re <= shift_reg_287_re;
    shift_reg_288_im <= shift_reg_287_im;
    shift_reg_289_re <= shift_reg_288_re;
    shift_reg_289_im <= shift_reg_288_im;
    shift_reg_290_re <= shift_reg_289_re;
    shift_reg_290_im <= shift_reg_289_im;
    shift_reg_291_re <= shift_reg_290_re;
    shift_reg_291_im <= shift_reg_290_im;
    shift_reg_292_re <= shift_reg_291_re;
    shift_reg_292_im <= shift_reg_291_im;
    shift_reg_293_re <= shift_reg_292_re;
    shift_reg_293_im <= shift_reg_292_im;
    shift_reg_294_re <= shift_reg_293_re;
    shift_reg_294_im <= shift_reg_293_im;
    shift_reg_295_re <= shift_reg_294_re;
    shift_reg_295_im <= shift_reg_294_im;
    shift_reg_296_re <= shift_reg_295_re;
    shift_reg_296_im <= shift_reg_295_im;
    shift_reg_297_re <= shift_reg_296_re;
    shift_reg_297_im <= shift_reg_296_im;
    shift_reg_298_re <= shift_reg_297_re;
    shift_reg_298_im <= shift_reg_297_im;
    shift_reg_299_re <= shift_reg_298_re;
    shift_reg_299_im <= shift_reg_298_im;
    shift_reg_300_re <= shift_reg_299_re;
    shift_reg_300_im <= shift_reg_299_im;
    shift_reg_301_re <= shift_reg_300_re;
    shift_reg_301_im <= shift_reg_300_im;
    shift_reg_302_re <= shift_reg_301_re;
    shift_reg_302_im <= shift_reg_301_im;
    shift_reg_303_re <= shift_reg_302_re;
    shift_reg_303_im <= shift_reg_302_im;
    shift_reg_304_re <= shift_reg_303_re;
    shift_reg_304_im <= shift_reg_303_im;
    shift_reg_305_re <= shift_reg_304_re;
    shift_reg_305_im <= shift_reg_304_im;
    shift_reg_306_re <= shift_reg_305_re;
    shift_reg_306_im <= shift_reg_305_im;
    shift_reg_307_re <= shift_reg_306_re;
    shift_reg_307_im <= shift_reg_306_im;
    shift_reg_308_re <= shift_reg_307_re;
    shift_reg_308_im <= shift_reg_307_im;
    shift_reg_309_re <= shift_reg_308_re;
    shift_reg_309_im <= shift_reg_308_im;
    shift_reg_310_re <= shift_reg_309_re;
    shift_reg_310_im <= shift_reg_309_im;
    shift_reg_311_re <= shift_reg_310_re;
    shift_reg_311_im <= shift_reg_310_im;
    shift_reg_312_re <= shift_reg_311_re;
    shift_reg_312_im <= shift_reg_311_im;
    shift_reg_313_re <= shift_reg_312_re;
    shift_reg_313_im <= shift_reg_312_im;
    shift_reg_314_re <= shift_reg_313_re;
    shift_reg_314_im <= shift_reg_313_im;
    shift_reg_315_re <= shift_reg_314_re;
    shift_reg_315_im <= shift_reg_314_im;
    shift_reg_316_re <= shift_reg_315_re;
    shift_reg_316_im <= shift_reg_315_im;
    shift_reg_317_re <= shift_reg_316_re;
    shift_reg_317_im <= shift_reg_316_im;
    shift_reg_318_re <= shift_reg_317_re;
    shift_reg_318_im <= shift_reg_317_im;
    shift_reg_319_re <= shift_reg_318_re;
    shift_reg_319_im <= shift_reg_318_im;
    shift_reg_320_re <= shift_reg_319_re;
    shift_reg_320_im <= shift_reg_319_im;
    shift_reg_321_re <= shift_reg_320_re;
    shift_reg_321_im <= shift_reg_320_im;
    shift_reg_322_re <= shift_reg_321_re;
    shift_reg_322_im <= shift_reg_321_im;
    shift_reg_323_re <= shift_reg_322_re;
    shift_reg_323_im <= shift_reg_322_im;
    shift_reg_324_re <= shift_reg_323_re;
    shift_reg_324_im <= shift_reg_323_im;
    shift_reg_325_re <= shift_reg_324_re;
    shift_reg_325_im <= shift_reg_324_im;
    shift_reg_326_re <= shift_reg_325_re;
    shift_reg_326_im <= shift_reg_325_im;
    shift_reg_327_re <= shift_reg_326_re;
    shift_reg_327_im <= shift_reg_326_im;
    shift_reg_328_re <= shift_reg_327_re;
    shift_reg_328_im <= shift_reg_327_im;
    shift_reg_329_re <= shift_reg_328_re;
    shift_reg_329_im <= shift_reg_328_im;
    shift_reg_330_re <= shift_reg_329_re;
    shift_reg_330_im <= shift_reg_329_im;
    shift_reg_331_re <= shift_reg_330_re;
    shift_reg_331_im <= shift_reg_330_im;
    shift_reg_332_re <= shift_reg_331_re;
    shift_reg_332_im <= shift_reg_331_im;
    shift_reg_333_re <= shift_reg_332_re;
    shift_reg_333_im <= shift_reg_332_im;
    shift_reg_334_re <= shift_reg_333_re;
    shift_reg_334_im <= shift_reg_333_im;
    shift_reg_335_re <= shift_reg_334_re;
    shift_reg_335_im <= shift_reg_334_im;
    shift_reg_336_re <= shift_reg_335_re;
    shift_reg_336_im <= shift_reg_335_im;
    shift_reg_337_re <= shift_reg_336_re;
    shift_reg_337_im <= shift_reg_336_im;
    shift_reg_338_re <= shift_reg_337_re;
    shift_reg_338_im <= shift_reg_337_im;
    shift_reg_339_re <= shift_reg_338_re;
    shift_reg_339_im <= shift_reg_338_im;
    shift_reg_340_re <= shift_reg_339_re;
    shift_reg_340_im <= shift_reg_339_im;
    shift_reg_341_re <= shift_reg_340_re;
    shift_reg_341_im <= shift_reg_340_im;
    shift_reg_342_re <= shift_reg_341_re;
    shift_reg_342_im <= shift_reg_341_im;
    shift_reg_343_re <= shift_reg_342_re;
    shift_reg_343_im <= shift_reg_342_im;
    shift_reg_344_re <= shift_reg_343_re;
    shift_reg_344_im <= shift_reg_343_im;
    shift_reg_345_re <= shift_reg_344_re;
    shift_reg_345_im <= shift_reg_344_im;
    shift_reg_346_re <= shift_reg_345_re;
    shift_reg_346_im <= shift_reg_345_im;
    shift_reg_347_re <= shift_reg_346_re;
    shift_reg_347_im <= shift_reg_346_im;
    shift_reg_348_re <= shift_reg_347_re;
    shift_reg_348_im <= shift_reg_347_im;
    shift_reg_349_re <= shift_reg_348_re;
    shift_reg_349_im <= shift_reg_348_im;
    shift_reg_350_re <= shift_reg_349_re;
    shift_reg_350_im <= shift_reg_349_im;
    shift_reg_351_re <= shift_reg_350_re;
    shift_reg_351_im <= shift_reg_350_im;
    shift_reg_352_re <= shift_reg_351_re;
    shift_reg_352_im <= shift_reg_351_im;
    shift_reg_353_re <= shift_reg_352_re;
    shift_reg_353_im <= shift_reg_352_im;
    shift_reg_354_re <= shift_reg_353_re;
    shift_reg_354_im <= shift_reg_353_im;
    shift_reg_355_re <= shift_reg_354_re;
    shift_reg_355_im <= shift_reg_354_im;
    shift_reg_356_re <= shift_reg_355_re;
    shift_reg_356_im <= shift_reg_355_im;
    shift_reg_357_re <= shift_reg_356_re;
    shift_reg_357_im <= shift_reg_356_im;
    shift_reg_358_re <= shift_reg_357_re;
    shift_reg_358_im <= shift_reg_357_im;
    shift_reg_359_re <= shift_reg_358_re;
    shift_reg_359_im <= shift_reg_358_im;
    shift_reg_360_re <= shift_reg_359_re;
    shift_reg_360_im <= shift_reg_359_im;
    shift_reg_361_re <= shift_reg_360_re;
    shift_reg_361_im <= shift_reg_360_im;
    shift_reg_362_re <= shift_reg_361_re;
    shift_reg_362_im <= shift_reg_361_im;
    shift_reg_363_re <= shift_reg_362_re;
    shift_reg_363_im <= shift_reg_362_im;
    shift_reg_364_re <= shift_reg_363_re;
    shift_reg_364_im <= shift_reg_363_im;
    shift_reg_365_re <= shift_reg_364_re;
    shift_reg_365_im <= shift_reg_364_im;
    shift_reg_366_re <= shift_reg_365_re;
    shift_reg_366_im <= shift_reg_365_im;
    shift_reg_367_re <= shift_reg_366_re;
    shift_reg_367_im <= shift_reg_366_im;
    shift_reg_368_re <= shift_reg_367_re;
    shift_reg_368_im <= shift_reg_367_im;
    shift_reg_369_re <= shift_reg_368_re;
    shift_reg_369_im <= shift_reg_368_im;
    shift_reg_370_re <= shift_reg_369_re;
    shift_reg_370_im <= shift_reg_369_im;
    shift_reg_371_re <= shift_reg_370_re;
    shift_reg_371_im <= shift_reg_370_im;
    shift_reg_372_re <= shift_reg_371_re;
    shift_reg_372_im <= shift_reg_371_im;
    shift_reg_373_re <= shift_reg_372_re;
    shift_reg_373_im <= shift_reg_372_im;
    shift_reg_374_re <= shift_reg_373_re;
    shift_reg_374_im <= shift_reg_373_im;
    shift_reg_375_re <= shift_reg_374_re;
    shift_reg_375_im <= shift_reg_374_im;
    shift_reg_376_re <= shift_reg_375_re;
    shift_reg_376_im <= shift_reg_375_im;
    shift_reg_377_re <= shift_reg_376_re;
    shift_reg_377_im <= shift_reg_376_im;
    shift_reg_378_re <= shift_reg_377_re;
    shift_reg_378_im <= shift_reg_377_im;
    shift_reg_379_re <= shift_reg_378_re;
    shift_reg_379_im <= shift_reg_378_im;
    shift_reg_380_re <= shift_reg_379_re;
    shift_reg_380_im <= shift_reg_379_im;
    shift_reg_381_re <= shift_reg_380_re;
    shift_reg_381_im <= shift_reg_380_im;
    shift_reg_382_re <= shift_reg_381_re;
    shift_reg_382_im <= shift_reg_381_im;
    shift_reg_383_re <= shift_reg_382_re;
    shift_reg_383_im <= shift_reg_382_im;
    shift_reg_384_re <= shift_reg_383_re;
    shift_reg_384_im <= shift_reg_383_im;
    shift_reg_385_re <= shift_reg_384_re;
    shift_reg_385_im <= shift_reg_384_im;
    shift_reg_386_re <= shift_reg_385_re;
    shift_reg_386_im <= shift_reg_385_im;
    shift_reg_387_re <= shift_reg_386_re;
    shift_reg_387_im <= shift_reg_386_im;
    shift_reg_388_re <= shift_reg_387_re;
    shift_reg_388_im <= shift_reg_387_im;
    shift_reg_389_re <= shift_reg_388_re;
    shift_reg_389_im <= shift_reg_388_im;
    shift_reg_390_re <= shift_reg_389_re;
    shift_reg_390_im <= shift_reg_389_im;
    shift_reg_391_re <= shift_reg_390_re;
    shift_reg_391_im <= shift_reg_390_im;
    shift_reg_392_re <= shift_reg_391_re;
    shift_reg_392_im <= shift_reg_391_im;
    shift_reg_393_re <= shift_reg_392_re;
    shift_reg_393_im <= shift_reg_392_im;
    shift_reg_394_re <= shift_reg_393_re;
    shift_reg_394_im <= shift_reg_393_im;
    shift_reg_395_re <= shift_reg_394_re;
    shift_reg_395_im <= shift_reg_394_im;
    shift_reg_396_re <= shift_reg_395_re;
    shift_reg_396_im <= shift_reg_395_im;
    shift_reg_397_re <= shift_reg_396_re;
    shift_reg_397_im <= shift_reg_396_im;
    shift_reg_398_re <= shift_reg_397_re;
    shift_reg_398_im <= shift_reg_397_im;
    shift_reg_399_re <= shift_reg_398_re;
    shift_reg_399_im <= shift_reg_398_im;
    shift_reg_400_re <= shift_reg_399_re;
    shift_reg_400_im <= shift_reg_399_im;
    shift_reg_401_re <= shift_reg_400_re;
    shift_reg_401_im <= shift_reg_400_im;
    shift_reg_402_re <= shift_reg_401_re;
    shift_reg_402_im <= shift_reg_401_im;
    shift_reg_403_re <= shift_reg_402_re;
    shift_reg_403_im <= shift_reg_402_im;
    shift_reg_404_re <= shift_reg_403_re;
    shift_reg_404_im <= shift_reg_403_im;
    shift_reg_405_re <= shift_reg_404_re;
    shift_reg_405_im <= shift_reg_404_im;
    shift_reg_406_re <= shift_reg_405_re;
    shift_reg_406_im <= shift_reg_405_im;
    shift_reg_407_re <= shift_reg_406_re;
    shift_reg_407_im <= shift_reg_406_im;
    shift_reg_408_re <= shift_reg_407_re;
    shift_reg_408_im <= shift_reg_407_im;
    shift_reg_409_re <= shift_reg_408_re;
    shift_reg_409_im <= shift_reg_408_im;
    shift_reg_410_re <= shift_reg_409_re;
    shift_reg_410_im <= shift_reg_409_im;
    shift_reg_411_re <= shift_reg_410_re;
    shift_reg_411_im <= shift_reg_410_im;
    shift_reg_412_re <= shift_reg_411_re;
    shift_reg_412_im <= shift_reg_411_im;
    shift_reg_413_re <= shift_reg_412_re;
    shift_reg_413_im <= shift_reg_412_im;
    shift_reg_414_re <= shift_reg_413_re;
    shift_reg_414_im <= shift_reg_413_im;
    shift_reg_415_re <= shift_reg_414_re;
    shift_reg_415_im <= shift_reg_414_im;
    shift_reg_416_re <= shift_reg_415_re;
    shift_reg_416_im <= shift_reg_415_im;
    shift_reg_417_re <= shift_reg_416_re;
    shift_reg_417_im <= shift_reg_416_im;
    shift_reg_418_re <= shift_reg_417_re;
    shift_reg_418_im <= shift_reg_417_im;
    shift_reg_419_re <= shift_reg_418_re;
    shift_reg_419_im <= shift_reg_418_im;
    shift_reg_420_re <= shift_reg_419_re;
    shift_reg_420_im <= shift_reg_419_im;
    shift_reg_421_re <= shift_reg_420_re;
    shift_reg_421_im <= shift_reg_420_im;
    shift_reg_422_re <= shift_reg_421_re;
    shift_reg_422_im <= shift_reg_421_im;
    shift_reg_423_re <= shift_reg_422_re;
    shift_reg_423_im <= shift_reg_422_im;
    shift_reg_424_re <= shift_reg_423_re;
    shift_reg_424_im <= shift_reg_423_im;
    shift_reg_425_re <= shift_reg_424_re;
    shift_reg_425_im <= shift_reg_424_im;
    shift_reg_426_re <= shift_reg_425_re;
    shift_reg_426_im <= shift_reg_425_im;
    shift_reg_427_re <= shift_reg_426_re;
    shift_reg_427_im <= shift_reg_426_im;
    shift_reg_428_re <= shift_reg_427_re;
    shift_reg_428_im <= shift_reg_427_im;
    shift_reg_429_re <= shift_reg_428_re;
    shift_reg_429_im <= shift_reg_428_im;
    shift_reg_430_re <= shift_reg_429_re;
    shift_reg_430_im <= shift_reg_429_im;
    shift_reg_431_re <= shift_reg_430_re;
    shift_reg_431_im <= shift_reg_430_im;
    shift_reg_432_re <= shift_reg_431_re;
    shift_reg_432_im <= shift_reg_431_im;
    shift_reg_433_re <= shift_reg_432_re;
    shift_reg_433_im <= shift_reg_432_im;
    shift_reg_434_re <= shift_reg_433_re;
    shift_reg_434_im <= shift_reg_433_im;
    shift_reg_435_re <= shift_reg_434_re;
    shift_reg_435_im <= shift_reg_434_im;
    shift_reg_436_re <= shift_reg_435_re;
    shift_reg_436_im <= shift_reg_435_im;
    shift_reg_437_re <= shift_reg_436_re;
    shift_reg_437_im <= shift_reg_436_im;
    shift_reg_438_re <= shift_reg_437_re;
    shift_reg_438_im <= shift_reg_437_im;
    shift_reg_439_re <= shift_reg_438_re;
    shift_reg_439_im <= shift_reg_438_im;
    shift_reg_440_re <= shift_reg_439_re;
    shift_reg_440_im <= shift_reg_439_im;
    shift_reg_441_re <= shift_reg_440_re;
    shift_reg_441_im <= shift_reg_440_im;
    shift_reg_442_re <= shift_reg_441_re;
    shift_reg_442_im <= shift_reg_441_im;
    shift_reg_443_re <= shift_reg_442_re;
    shift_reg_443_im <= shift_reg_442_im;
    shift_reg_444_re <= shift_reg_443_re;
    shift_reg_444_im <= shift_reg_443_im;
    shift_reg_445_re <= shift_reg_444_re;
    shift_reg_445_im <= shift_reg_444_im;
    shift_reg_446_re <= shift_reg_445_re;
    shift_reg_446_im <= shift_reg_445_im;
    shift_reg_447_re <= shift_reg_446_re;
    shift_reg_447_im <= shift_reg_446_im;
    shift_reg_448_re <= shift_reg_447_re;
    shift_reg_448_im <= shift_reg_447_im;
    shift_reg_449_re <= shift_reg_448_re;
    shift_reg_449_im <= shift_reg_448_im;
    shift_reg_450_re <= shift_reg_449_re;
    shift_reg_450_im <= shift_reg_449_im;
    shift_reg_451_re <= shift_reg_450_re;
    shift_reg_451_im <= shift_reg_450_im;
    shift_reg_452_re <= shift_reg_451_re;
    shift_reg_452_im <= shift_reg_451_im;
    shift_reg_453_re <= shift_reg_452_re;
    shift_reg_453_im <= shift_reg_452_im;
    shift_reg_454_re <= shift_reg_453_re;
    shift_reg_454_im <= shift_reg_453_im;
    shift_reg_455_re <= shift_reg_454_re;
    shift_reg_455_im <= shift_reg_454_im;
    shift_reg_456_re <= shift_reg_455_re;
    shift_reg_456_im <= shift_reg_455_im;
    shift_reg_457_re <= shift_reg_456_re;
    shift_reg_457_im <= shift_reg_456_im;
    shift_reg_458_re <= shift_reg_457_re;
    shift_reg_458_im <= shift_reg_457_im;
    shift_reg_459_re <= shift_reg_458_re;
    shift_reg_459_im <= shift_reg_458_im;
    shift_reg_460_re <= shift_reg_459_re;
    shift_reg_460_im <= shift_reg_459_im;
    shift_reg_461_re <= shift_reg_460_re;
    shift_reg_461_im <= shift_reg_460_im;
    shift_reg_462_re <= shift_reg_461_re;
    shift_reg_462_im <= shift_reg_461_im;
    shift_reg_463_re <= shift_reg_462_re;
    shift_reg_463_im <= shift_reg_462_im;
    shift_reg_464_re <= shift_reg_463_re;
    shift_reg_464_im <= shift_reg_463_im;
    shift_reg_465_re <= shift_reg_464_re;
    shift_reg_465_im <= shift_reg_464_im;
    shift_reg_466_re <= shift_reg_465_re;
    shift_reg_466_im <= shift_reg_465_im;
    shift_reg_467_re <= shift_reg_466_re;
    shift_reg_467_im <= shift_reg_466_im;
    shift_reg_468_re <= shift_reg_467_re;
    shift_reg_468_im <= shift_reg_467_im;
    shift_reg_469_re <= shift_reg_468_re;
    shift_reg_469_im <= shift_reg_468_im;
    shift_reg_470_re <= shift_reg_469_re;
    shift_reg_470_im <= shift_reg_469_im;
    shift_reg_471_re <= shift_reg_470_re;
    shift_reg_471_im <= shift_reg_470_im;
    shift_reg_472_re <= shift_reg_471_re;
    shift_reg_472_im <= shift_reg_471_im;
    shift_reg_473_re <= shift_reg_472_re;
    shift_reg_473_im <= shift_reg_472_im;
    shift_reg_474_re <= shift_reg_473_re;
    shift_reg_474_im <= shift_reg_473_im;
    shift_reg_475_re <= shift_reg_474_re;
    shift_reg_475_im <= shift_reg_474_im;
    shift_reg_476_re <= shift_reg_475_re;
    shift_reg_476_im <= shift_reg_475_im;
    shift_reg_477_re <= shift_reg_476_re;
    shift_reg_477_im <= shift_reg_476_im;
    shift_reg_478_re <= shift_reg_477_re;
    shift_reg_478_im <= shift_reg_477_im;
    shift_reg_479_re <= shift_reg_478_re;
    shift_reg_479_im <= shift_reg_478_im;
    shift_reg_480_re <= shift_reg_479_re;
    shift_reg_480_im <= shift_reg_479_im;
    shift_reg_481_re <= shift_reg_480_re;
    shift_reg_481_im <= shift_reg_480_im;
    shift_reg_482_re <= shift_reg_481_re;
    shift_reg_482_im <= shift_reg_481_im;
    shift_reg_483_re <= shift_reg_482_re;
    shift_reg_483_im <= shift_reg_482_im;
    shift_reg_484_re <= shift_reg_483_re;
    shift_reg_484_im <= shift_reg_483_im;
    shift_reg_485_re <= shift_reg_484_re;
    shift_reg_485_im <= shift_reg_484_im;
    shift_reg_486_re <= shift_reg_485_re;
    shift_reg_486_im <= shift_reg_485_im;
    shift_reg_487_re <= shift_reg_486_re;
    shift_reg_487_im <= shift_reg_486_im;
    shift_reg_488_re <= shift_reg_487_re;
    shift_reg_488_im <= shift_reg_487_im;
    shift_reg_489_re <= shift_reg_488_re;
    shift_reg_489_im <= shift_reg_488_im;
    shift_reg_490_re <= shift_reg_489_re;
    shift_reg_490_im <= shift_reg_489_im;
    shift_reg_491_re <= shift_reg_490_re;
    shift_reg_491_im <= shift_reg_490_im;
    shift_reg_492_re <= shift_reg_491_re;
    shift_reg_492_im <= shift_reg_491_im;
    shift_reg_493_re <= shift_reg_492_re;
    shift_reg_493_im <= shift_reg_492_im;
    shift_reg_494_re <= shift_reg_493_re;
    shift_reg_494_im <= shift_reg_493_im;
    shift_reg_495_re <= shift_reg_494_re;
    shift_reg_495_im <= shift_reg_494_im;
    shift_reg_496_re <= shift_reg_495_re;
    shift_reg_496_im <= shift_reg_495_im;
    shift_reg_497_re <= shift_reg_496_re;
    shift_reg_497_im <= shift_reg_496_im;
    shift_reg_498_re <= shift_reg_497_re;
    shift_reg_498_im <= shift_reg_497_im;
    shift_reg_499_re <= shift_reg_498_re;
    shift_reg_499_im <= shift_reg_498_im;
    shift_reg_500_re <= shift_reg_499_re;
    shift_reg_500_im <= shift_reg_499_im;
    shift_reg_501_re <= shift_reg_500_re;
    shift_reg_501_im <= shift_reg_500_im;
    shift_reg_502_re <= shift_reg_501_re;
    shift_reg_502_im <= shift_reg_501_im;
    shift_reg_503_re <= shift_reg_502_re;
    shift_reg_503_im <= shift_reg_502_im;
    shift_reg_504_re <= shift_reg_503_re;
    shift_reg_504_im <= shift_reg_503_im;
    shift_reg_505_re <= shift_reg_504_re;
    shift_reg_505_im <= shift_reg_504_im;
    shift_reg_506_re <= shift_reg_505_re;
    shift_reg_506_im <= shift_reg_505_im;
    shift_reg_507_re <= shift_reg_506_re;
    shift_reg_507_im <= shift_reg_506_im;
    shift_reg_508_re <= shift_reg_507_re;
    shift_reg_508_im <= shift_reg_507_im;
    shift_reg_509_re <= shift_reg_508_re;
    shift_reg_509_im <= shift_reg_508_im;
    shift_reg_510_re <= shift_reg_509_re;
    shift_reg_510_im <= shift_reg_509_im;
    shift_reg_511_re <= shift_reg_510_re;
    shift_reg_511_im <= shift_reg_510_im;
    shift_reg_512_re <= shift_reg_511_re;
    shift_reg_512_im <= shift_reg_511_im;
    shift_reg_513_re <= shift_reg_512_re;
    shift_reg_513_im <= shift_reg_512_im;
    shift_reg_514_re <= shift_reg_513_re;
    shift_reg_514_im <= shift_reg_513_im;
    shift_reg_515_re <= shift_reg_514_re;
    shift_reg_515_im <= shift_reg_514_im;
    shift_reg_516_re <= shift_reg_515_re;
    shift_reg_516_im <= shift_reg_515_im;
    shift_reg_517_re <= shift_reg_516_re;
    shift_reg_517_im <= shift_reg_516_im;
    shift_reg_518_re <= shift_reg_517_re;
    shift_reg_518_im <= shift_reg_517_im;
    shift_reg_519_re <= shift_reg_518_re;
    shift_reg_519_im <= shift_reg_518_im;
    shift_reg_520_re <= shift_reg_519_re;
    shift_reg_520_im <= shift_reg_519_im;
    shift_reg_521_re <= shift_reg_520_re;
    shift_reg_521_im <= shift_reg_520_im;
    shift_reg_522_re <= shift_reg_521_re;
    shift_reg_522_im <= shift_reg_521_im;
    shift_reg_523_re <= shift_reg_522_re;
    shift_reg_523_im <= shift_reg_522_im;
    shift_reg_524_re <= shift_reg_523_re;
    shift_reg_524_im <= shift_reg_523_im;
    shift_reg_525_re <= shift_reg_524_re;
    shift_reg_525_im <= shift_reg_524_im;
    shift_reg_526_re <= shift_reg_525_re;
    shift_reg_526_im <= shift_reg_525_im;
    shift_reg_527_re <= shift_reg_526_re;
    shift_reg_527_im <= shift_reg_526_im;
    shift_reg_528_re <= shift_reg_527_re;
    shift_reg_528_im <= shift_reg_527_im;
    shift_reg_529_re <= shift_reg_528_re;
    shift_reg_529_im <= shift_reg_528_im;
    shift_reg_530_re <= shift_reg_529_re;
    shift_reg_530_im <= shift_reg_529_im;
    shift_reg_531_re <= shift_reg_530_re;
    shift_reg_531_im <= shift_reg_530_im;
    shift_reg_532_re <= shift_reg_531_re;
    shift_reg_532_im <= shift_reg_531_im;
    shift_reg_533_re <= shift_reg_532_re;
    shift_reg_533_im <= shift_reg_532_im;
    shift_reg_534_re <= shift_reg_533_re;
    shift_reg_534_im <= shift_reg_533_im;
    shift_reg_535_re <= shift_reg_534_re;
    shift_reg_535_im <= shift_reg_534_im;
    shift_reg_536_re <= shift_reg_535_re;
    shift_reg_536_im <= shift_reg_535_im;
    shift_reg_537_re <= shift_reg_536_re;
    shift_reg_537_im <= shift_reg_536_im;
    shift_reg_538_re <= shift_reg_537_re;
    shift_reg_538_im <= shift_reg_537_im;
    shift_reg_539_re <= shift_reg_538_re;
    shift_reg_539_im <= shift_reg_538_im;
    shift_reg_540_re <= shift_reg_539_re;
    shift_reg_540_im <= shift_reg_539_im;
    shift_reg_541_re <= shift_reg_540_re;
    shift_reg_541_im <= shift_reg_540_im;
    shift_reg_542_re <= shift_reg_541_re;
    shift_reg_542_im <= shift_reg_541_im;
    shift_reg_543_re <= shift_reg_542_re;
    shift_reg_543_im <= shift_reg_542_im;
    shift_reg_544_re <= shift_reg_543_re;
    shift_reg_544_im <= shift_reg_543_im;
    shift_reg_545_re <= shift_reg_544_re;
    shift_reg_545_im <= shift_reg_544_im;
    shift_reg_546_re <= shift_reg_545_re;
    shift_reg_546_im <= shift_reg_545_im;
    shift_reg_547_re <= shift_reg_546_re;
    shift_reg_547_im <= shift_reg_546_im;
    shift_reg_548_re <= shift_reg_547_re;
    shift_reg_548_im <= shift_reg_547_im;
    shift_reg_549_re <= shift_reg_548_re;
    shift_reg_549_im <= shift_reg_548_im;
    shift_reg_550_re <= shift_reg_549_re;
    shift_reg_550_im <= shift_reg_549_im;
    shift_reg_551_re <= shift_reg_550_re;
    shift_reg_551_im <= shift_reg_550_im;
    shift_reg_552_re <= shift_reg_551_re;
    shift_reg_552_im <= shift_reg_551_im;
    shift_reg_553_re <= shift_reg_552_re;
    shift_reg_553_im <= shift_reg_552_im;
    shift_reg_554_re <= shift_reg_553_re;
    shift_reg_554_im <= shift_reg_553_im;
    shift_reg_555_re <= shift_reg_554_re;
    shift_reg_555_im <= shift_reg_554_im;
    shift_reg_556_re <= shift_reg_555_re;
    shift_reg_556_im <= shift_reg_555_im;
    shift_reg_557_re <= shift_reg_556_re;
    shift_reg_557_im <= shift_reg_556_im;
    shift_reg_558_re <= shift_reg_557_re;
    shift_reg_558_im <= shift_reg_557_im;
    shift_reg_559_re <= shift_reg_558_re;
    shift_reg_559_im <= shift_reg_558_im;
    shift_reg_560_re <= shift_reg_559_re;
    shift_reg_560_im <= shift_reg_559_im;
    shift_reg_561_re <= shift_reg_560_re;
    shift_reg_561_im <= shift_reg_560_im;
    shift_reg_562_re <= shift_reg_561_re;
    shift_reg_562_im <= shift_reg_561_im;
    shift_reg_563_re <= shift_reg_562_re;
    shift_reg_563_im <= shift_reg_562_im;
    shift_reg_564_re <= shift_reg_563_re;
    shift_reg_564_im <= shift_reg_563_im;
    shift_reg_565_re <= shift_reg_564_re;
    shift_reg_565_im <= shift_reg_564_im;
    shift_reg_566_re <= shift_reg_565_re;
    shift_reg_566_im <= shift_reg_565_im;
    shift_reg_567_re <= shift_reg_566_re;
    shift_reg_567_im <= shift_reg_566_im;
    shift_reg_568_re <= shift_reg_567_re;
    shift_reg_568_im <= shift_reg_567_im;
    shift_reg_569_re <= shift_reg_568_re;
    shift_reg_569_im <= shift_reg_568_im;
    shift_reg_570_re <= shift_reg_569_re;
    shift_reg_570_im <= shift_reg_569_im;
    shift_reg_571_re <= shift_reg_570_re;
    shift_reg_571_im <= shift_reg_570_im;
    shift_reg_572_re <= shift_reg_571_re;
    shift_reg_572_im <= shift_reg_571_im;
    shift_reg_573_re <= shift_reg_572_re;
    shift_reg_573_im <= shift_reg_572_im;
    shift_reg_574_re <= shift_reg_573_re;
    shift_reg_574_im <= shift_reg_573_im;
    shift_reg_575_re <= shift_reg_574_re;
    shift_reg_575_im <= shift_reg_574_im;
    shift_reg_576_re <= shift_reg_575_re;
    shift_reg_576_im <= shift_reg_575_im;
    shift_reg_577_re <= shift_reg_576_re;
    shift_reg_577_im <= shift_reg_576_im;
    shift_reg_578_re <= shift_reg_577_re;
    shift_reg_578_im <= shift_reg_577_im;
    shift_reg_579_re <= shift_reg_578_re;
    shift_reg_579_im <= shift_reg_578_im;
    shift_reg_580_re <= shift_reg_579_re;
    shift_reg_580_im <= shift_reg_579_im;
    shift_reg_581_re <= shift_reg_580_re;
    shift_reg_581_im <= shift_reg_580_im;
    shift_reg_582_re <= shift_reg_581_re;
    shift_reg_582_im <= shift_reg_581_im;
    shift_reg_583_re <= shift_reg_582_re;
    shift_reg_583_im <= shift_reg_582_im;
    shift_reg_584_re <= shift_reg_583_re;
    shift_reg_584_im <= shift_reg_583_im;
    shift_reg_585_re <= shift_reg_584_re;
    shift_reg_585_im <= shift_reg_584_im;
    shift_reg_586_re <= shift_reg_585_re;
    shift_reg_586_im <= shift_reg_585_im;
    shift_reg_587_re <= shift_reg_586_re;
    shift_reg_587_im <= shift_reg_586_im;
    shift_reg_588_re <= shift_reg_587_re;
    shift_reg_588_im <= shift_reg_587_im;
    shift_reg_589_re <= shift_reg_588_re;
    shift_reg_589_im <= shift_reg_588_im;
    shift_reg_590_re <= shift_reg_589_re;
    shift_reg_590_im <= shift_reg_589_im;
    shift_reg_591_re <= shift_reg_590_re;
    shift_reg_591_im <= shift_reg_590_im;
    shift_reg_592_re <= shift_reg_591_re;
    shift_reg_592_im <= shift_reg_591_im;
    shift_reg_593_re <= shift_reg_592_re;
    shift_reg_593_im <= shift_reg_592_im;
    shift_reg_594_re <= shift_reg_593_re;
    shift_reg_594_im <= shift_reg_593_im;
    shift_reg_595_re <= shift_reg_594_re;
    shift_reg_595_im <= shift_reg_594_im;
    shift_reg_596_re <= shift_reg_595_re;
    shift_reg_596_im <= shift_reg_595_im;
    shift_reg_597_re <= shift_reg_596_re;
    shift_reg_597_im <= shift_reg_596_im;
    shift_reg_598_re <= shift_reg_597_re;
    shift_reg_598_im <= shift_reg_597_im;
    shift_reg_599_re <= shift_reg_598_re;
    shift_reg_599_im <= shift_reg_598_im;
    shift_reg_600_re <= shift_reg_599_re;
    shift_reg_600_im <= shift_reg_599_im;
    shift_reg_601_re <= shift_reg_600_re;
    shift_reg_601_im <= shift_reg_600_im;
    shift_reg_602_re <= shift_reg_601_re;
    shift_reg_602_im <= shift_reg_601_im;
    shift_reg_603_re <= shift_reg_602_re;
    shift_reg_603_im <= shift_reg_602_im;
    shift_reg_604_re <= shift_reg_603_re;
    shift_reg_604_im <= shift_reg_603_im;
    shift_reg_605_re <= shift_reg_604_re;
    shift_reg_605_im <= shift_reg_604_im;
    shift_reg_606_re <= shift_reg_605_re;
    shift_reg_606_im <= shift_reg_605_im;
    shift_reg_607_re <= shift_reg_606_re;
    shift_reg_607_im <= shift_reg_606_im;
    shift_reg_608_re <= shift_reg_607_re;
    shift_reg_608_im <= shift_reg_607_im;
    shift_reg_609_re <= shift_reg_608_re;
    shift_reg_609_im <= shift_reg_608_im;
    shift_reg_610_re <= shift_reg_609_re;
    shift_reg_610_im <= shift_reg_609_im;
    shift_reg_611_re <= shift_reg_610_re;
    shift_reg_611_im <= shift_reg_610_im;
    shift_reg_612_re <= shift_reg_611_re;
    shift_reg_612_im <= shift_reg_611_im;
    shift_reg_613_re <= shift_reg_612_re;
    shift_reg_613_im <= shift_reg_612_im;
    shift_reg_614_re <= shift_reg_613_re;
    shift_reg_614_im <= shift_reg_613_im;
    shift_reg_615_re <= shift_reg_614_re;
    shift_reg_615_im <= shift_reg_614_im;
    shift_reg_616_re <= shift_reg_615_re;
    shift_reg_616_im <= shift_reg_615_im;
    shift_reg_617_re <= shift_reg_616_re;
    shift_reg_617_im <= shift_reg_616_im;
    shift_reg_618_re <= shift_reg_617_re;
    shift_reg_618_im <= shift_reg_617_im;
    shift_reg_619_re <= shift_reg_618_re;
    shift_reg_619_im <= shift_reg_618_im;
    shift_reg_620_re <= shift_reg_619_re;
    shift_reg_620_im <= shift_reg_619_im;
    shift_reg_621_re <= shift_reg_620_re;
    shift_reg_621_im <= shift_reg_620_im;
    shift_reg_622_re <= shift_reg_621_re;
    shift_reg_622_im <= shift_reg_621_im;
    shift_reg_623_re <= shift_reg_622_re;
    shift_reg_623_im <= shift_reg_622_im;
    shift_reg_624_re <= shift_reg_623_re;
    shift_reg_624_im <= shift_reg_623_im;
    shift_reg_625_re <= shift_reg_624_re;
    shift_reg_625_im <= shift_reg_624_im;
    shift_reg_626_re <= shift_reg_625_re;
    shift_reg_626_im <= shift_reg_625_im;
    shift_reg_627_re <= shift_reg_626_re;
    shift_reg_627_im <= shift_reg_626_im;
    shift_reg_628_re <= shift_reg_627_re;
    shift_reg_628_im <= shift_reg_627_im;
    shift_reg_629_re <= shift_reg_628_re;
    shift_reg_629_im <= shift_reg_628_im;
    shift_reg_630_re <= shift_reg_629_re;
    shift_reg_630_im <= shift_reg_629_im;
    shift_reg_631_re <= shift_reg_630_re;
    shift_reg_631_im <= shift_reg_630_im;
    shift_reg_632_re <= shift_reg_631_re;
    shift_reg_632_im <= shift_reg_631_im;
    shift_reg_633_re <= shift_reg_632_re;
    shift_reg_633_im <= shift_reg_632_im;
    shift_reg_634_re <= shift_reg_633_re;
    shift_reg_634_im <= shift_reg_633_im;
    shift_reg_635_re <= shift_reg_634_re;
    shift_reg_635_im <= shift_reg_634_im;
    shift_reg_636_re <= shift_reg_635_re;
    shift_reg_636_im <= shift_reg_635_im;
    shift_reg_637_re <= shift_reg_636_re;
    shift_reg_637_im <= shift_reg_636_im;
    shift_reg_638_re <= shift_reg_637_re;
    shift_reg_638_im <= shift_reg_637_im;
    shift_reg_639_re <= shift_reg_638_re;
    shift_reg_639_im <= shift_reg_638_im;
    shift_reg_640_re <= shift_reg_639_re;
    shift_reg_640_im <= shift_reg_639_im;
    shift_reg_641_re <= shift_reg_640_re;
    shift_reg_641_im <= shift_reg_640_im;
    shift_reg_642_re <= shift_reg_641_re;
    shift_reg_642_im <= shift_reg_641_im;
    shift_reg_643_re <= shift_reg_642_re;
    shift_reg_643_im <= shift_reg_642_im;
    shift_reg_644_re <= shift_reg_643_re;
    shift_reg_644_im <= shift_reg_643_im;
    shift_reg_645_re <= shift_reg_644_re;
    shift_reg_645_im <= shift_reg_644_im;
    shift_reg_646_re <= shift_reg_645_re;
    shift_reg_646_im <= shift_reg_645_im;
    shift_reg_647_re <= shift_reg_646_re;
    shift_reg_647_im <= shift_reg_646_im;
    shift_reg_648_re <= shift_reg_647_re;
    shift_reg_648_im <= shift_reg_647_im;
    shift_reg_649_re <= shift_reg_648_re;
    shift_reg_649_im <= shift_reg_648_im;
    shift_reg_650_re <= shift_reg_649_re;
    shift_reg_650_im <= shift_reg_649_im;
    shift_reg_651_re <= shift_reg_650_re;
    shift_reg_651_im <= shift_reg_650_im;
    shift_reg_652_re <= shift_reg_651_re;
    shift_reg_652_im <= shift_reg_651_im;
    shift_reg_653_re <= shift_reg_652_re;
    shift_reg_653_im <= shift_reg_652_im;
    shift_reg_654_re <= shift_reg_653_re;
    shift_reg_654_im <= shift_reg_653_im;
    shift_reg_655_re <= shift_reg_654_re;
    shift_reg_655_im <= shift_reg_654_im;
    shift_reg_656_re <= shift_reg_655_re;
    shift_reg_656_im <= shift_reg_655_im;
    shift_reg_657_re <= shift_reg_656_re;
    shift_reg_657_im <= shift_reg_656_im;
    shift_reg_658_re <= shift_reg_657_re;
    shift_reg_658_im <= shift_reg_657_im;
    shift_reg_659_re <= shift_reg_658_re;
    shift_reg_659_im <= shift_reg_658_im;
    shift_reg_660_re <= shift_reg_659_re;
    shift_reg_660_im <= shift_reg_659_im;
    shift_reg_661_re <= shift_reg_660_re;
    shift_reg_661_im <= shift_reg_660_im;
    shift_reg_662_re <= shift_reg_661_re;
    shift_reg_662_im <= shift_reg_661_im;
    shift_reg_663_re <= shift_reg_662_re;
    shift_reg_663_im <= shift_reg_662_im;
    shift_reg_664_re <= shift_reg_663_re;
    shift_reg_664_im <= shift_reg_663_im;
    shift_reg_665_re <= shift_reg_664_re;
    shift_reg_665_im <= shift_reg_664_im;
    shift_reg_666_re <= shift_reg_665_re;
    shift_reg_666_im <= shift_reg_665_im;
    shift_reg_667_re <= shift_reg_666_re;
    shift_reg_667_im <= shift_reg_666_im;
    shift_reg_668_re <= shift_reg_667_re;
    shift_reg_668_im <= shift_reg_667_im;
    shift_reg_669_re <= shift_reg_668_re;
    shift_reg_669_im <= shift_reg_668_im;
    shift_reg_670_re <= shift_reg_669_re;
    shift_reg_670_im <= shift_reg_669_im;
    shift_reg_671_re <= shift_reg_670_re;
    shift_reg_671_im <= shift_reg_670_im;
    shift_reg_672_re <= shift_reg_671_re;
    shift_reg_672_im <= shift_reg_671_im;
    shift_reg_673_re <= shift_reg_672_re;
    shift_reg_673_im <= shift_reg_672_im;
    shift_reg_674_re <= shift_reg_673_re;
    shift_reg_674_im <= shift_reg_673_im;
    shift_reg_675_re <= shift_reg_674_re;
    shift_reg_675_im <= shift_reg_674_im;
    shift_reg_676_re <= shift_reg_675_re;
    shift_reg_676_im <= shift_reg_675_im;
    shift_reg_677_re <= shift_reg_676_re;
    shift_reg_677_im <= shift_reg_676_im;
    shift_reg_678_re <= shift_reg_677_re;
    shift_reg_678_im <= shift_reg_677_im;
    shift_reg_679_re <= shift_reg_678_re;
    shift_reg_679_im <= shift_reg_678_im;
    shift_reg_680_re <= shift_reg_679_re;
    shift_reg_680_im <= shift_reg_679_im;
    shift_reg_681_re <= shift_reg_680_re;
    shift_reg_681_im <= shift_reg_680_im;
    shift_reg_682_re <= shift_reg_681_re;
    shift_reg_682_im <= shift_reg_681_im;
    shift_reg_683_re <= shift_reg_682_re;
    shift_reg_683_im <= shift_reg_682_im;
    shift_reg_684_re <= shift_reg_683_re;
    shift_reg_684_im <= shift_reg_683_im;
    shift_reg_685_re <= shift_reg_684_re;
    shift_reg_685_im <= shift_reg_684_im;
    shift_reg_686_re <= shift_reg_685_re;
    shift_reg_686_im <= shift_reg_685_im;
    shift_reg_687_re <= shift_reg_686_re;
    shift_reg_687_im <= shift_reg_686_im;
    shift_reg_688_re <= shift_reg_687_re;
    shift_reg_688_im <= shift_reg_687_im;
    shift_reg_689_re <= shift_reg_688_re;
    shift_reg_689_im <= shift_reg_688_im;
    shift_reg_690_re <= shift_reg_689_re;
    shift_reg_690_im <= shift_reg_689_im;
    shift_reg_691_re <= shift_reg_690_re;
    shift_reg_691_im <= shift_reg_690_im;
    shift_reg_692_re <= shift_reg_691_re;
    shift_reg_692_im <= shift_reg_691_im;
    shift_reg_693_re <= shift_reg_692_re;
    shift_reg_693_im <= shift_reg_692_im;
    shift_reg_694_re <= shift_reg_693_re;
    shift_reg_694_im <= shift_reg_693_im;
    shift_reg_695_re <= shift_reg_694_re;
    shift_reg_695_im <= shift_reg_694_im;
    shift_reg_696_re <= shift_reg_695_re;
    shift_reg_696_im <= shift_reg_695_im;
    shift_reg_697_re <= shift_reg_696_re;
    shift_reg_697_im <= shift_reg_696_im;
    shift_reg_698_re <= shift_reg_697_re;
    shift_reg_698_im <= shift_reg_697_im;
    shift_reg_699_re <= shift_reg_698_re;
    shift_reg_699_im <= shift_reg_698_im;
    shift_reg_700_re <= shift_reg_699_re;
    shift_reg_700_im <= shift_reg_699_im;
    shift_reg_701_re <= shift_reg_700_re;
    shift_reg_701_im <= shift_reg_700_im;
    shift_reg_702_re <= shift_reg_701_re;
    shift_reg_702_im <= shift_reg_701_im;
    shift_reg_703_re <= shift_reg_702_re;
    shift_reg_703_im <= shift_reg_702_im;
    shift_reg_704_re <= shift_reg_703_re;
    shift_reg_704_im <= shift_reg_703_im;
    shift_reg_705_re <= shift_reg_704_re;
    shift_reg_705_im <= shift_reg_704_im;
    shift_reg_706_re <= shift_reg_705_re;
    shift_reg_706_im <= shift_reg_705_im;
    shift_reg_707_re <= shift_reg_706_re;
    shift_reg_707_im <= shift_reg_706_im;
    shift_reg_708_re <= shift_reg_707_re;
    shift_reg_708_im <= shift_reg_707_im;
    shift_reg_709_re <= shift_reg_708_re;
    shift_reg_709_im <= shift_reg_708_im;
    shift_reg_710_re <= shift_reg_709_re;
    shift_reg_710_im <= shift_reg_709_im;
    shift_reg_711_re <= shift_reg_710_re;
    shift_reg_711_im <= shift_reg_710_im;
    shift_reg_712_re <= shift_reg_711_re;
    shift_reg_712_im <= shift_reg_711_im;
    shift_reg_713_re <= shift_reg_712_re;
    shift_reg_713_im <= shift_reg_712_im;
    shift_reg_714_re <= shift_reg_713_re;
    shift_reg_714_im <= shift_reg_713_im;
    shift_reg_715_re <= shift_reg_714_re;
    shift_reg_715_im <= shift_reg_714_im;
    shift_reg_716_re <= shift_reg_715_re;
    shift_reg_716_im <= shift_reg_715_im;
    shift_reg_717_re <= shift_reg_716_re;
    shift_reg_717_im <= shift_reg_716_im;
    shift_reg_718_re <= shift_reg_717_re;
    shift_reg_718_im <= shift_reg_717_im;
    shift_reg_719_re <= shift_reg_718_re;
    shift_reg_719_im <= shift_reg_718_im;
    shift_reg_720_re <= shift_reg_719_re;
    shift_reg_720_im <= shift_reg_719_im;
    shift_reg_721_re <= shift_reg_720_re;
    shift_reg_721_im <= shift_reg_720_im;
    shift_reg_722_re <= shift_reg_721_re;
    shift_reg_722_im <= shift_reg_721_im;
    shift_reg_723_re <= shift_reg_722_re;
    shift_reg_723_im <= shift_reg_722_im;
    shift_reg_724_re <= shift_reg_723_re;
    shift_reg_724_im <= shift_reg_723_im;
    shift_reg_725_re <= shift_reg_724_re;
    shift_reg_725_im <= shift_reg_724_im;
    shift_reg_726_re <= shift_reg_725_re;
    shift_reg_726_im <= shift_reg_725_im;
    shift_reg_727_re <= shift_reg_726_re;
    shift_reg_727_im <= shift_reg_726_im;
    shift_reg_728_re <= shift_reg_727_re;
    shift_reg_728_im <= shift_reg_727_im;
    shift_reg_729_re <= shift_reg_728_re;
    shift_reg_729_im <= shift_reg_728_im;
    shift_reg_730_re <= shift_reg_729_re;
    shift_reg_730_im <= shift_reg_729_im;
    shift_reg_731_re <= shift_reg_730_re;
    shift_reg_731_im <= shift_reg_730_im;
    shift_reg_732_re <= shift_reg_731_re;
    shift_reg_732_im <= shift_reg_731_im;
    shift_reg_733_re <= shift_reg_732_re;
    shift_reg_733_im <= shift_reg_732_im;
    shift_reg_734_re <= shift_reg_733_re;
    shift_reg_734_im <= shift_reg_733_im;
    shift_reg_735_re <= shift_reg_734_re;
    shift_reg_735_im <= shift_reg_734_im;
    shift_reg_736_re <= shift_reg_735_re;
    shift_reg_736_im <= shift_reg_735_im;
    shift_reg_737_re <= shift_reg_736_re;
    shift_reg_737_im <= shift_reg_736_im;
    shift_reg_738_re <= shift_reg_737_re;
    shift_reg_738_im <= shift_reg_737_im;
    shift_reg_739_re <= shift_reg_738_re;
    shift_reg_739_im <= shift_reg_738_im;
    shift_reg_740_re <= shift_reg_739_re;
    shift_reg_740_im <= shift_reg_739_im;
    shift_reg_741_re <= shift_reg_740_re;
    shift_reg_741_im <= shift_reg_740_im;
    shift_reg_742_re <= shift_reg_741_re;
    shift_reg_742_im <= shift_reg_741_im;
    shift_reg_743_re <= shift_reg_742_re;
    shift_reg_743_im <= shift_reg_742_im;
    shift_reg_744_re <= shift_reg_743_re;
    shift_reg_744_im <= shift_reg_743_im;
    shift_reg_745_re <= shift_reg_744_re;
    shift_reg_745_im <= shift_reg_744_im;
    shift_reg_746_re <= shift_reg_745_re;
    shift_reg_746_im <= shift_reg_745_im;
    shift_reg_747_re <= shift_reg_746_re;
    shift_reg_747_im <= shift_reg_746_im;
    shift_reg_748_re <= shift_reg_747_re;
    shift_reg_748_im <= shift_reg_747_im;
    shift_reg_749_re <= shift_reg_748_re;
    shift_reg_749_im <= shift_reg_748_im;
    shift_reg_750_re <= shift_reg_749_re;
    shift_reg_750_im <= shift_reg_749_im;
    shift_reg_751_re <= shift_reg_750_re;
    shift_reg_751_im <= shift_reg_750_im;
    shift_reg_752_re <= shift_reg_751_re;
    shift_reg_752_im <= shift_reg_751_im;
    shift_reg_753_re <= shift_reg_752_re;
    shift_reg_753_im <= shift_reg_752_im;
    shift_reg_754_re <= shift_reg_753_re;
    shift_reg_754_im <= shift_reg_753_im;
    shift_reg_755_re <= shift_reg_754_re;
    shift_reg_755_im <= shift_reg_754_im;
    shift_reg_756_re <= shift_reg_755_re;
    shift_reg_756_im <= shift_reg_755_im;
    shift_reg_757_re <= shift_reg_756_re;
    shift_reg_757_im <= shift_reg_756_im;
    shift_reg_758_re <= shift_reg_757_re;
    shift_reg_758_im <= shift_reg_757_im;
    shift_reg_759_re <= shift_reg_758_re;
    shift_reg_759_im <= shift_reg_758_im;
    shift_reg_760_re <= shift_reg_759_re;
    shift_reg_760_im <= shift_reg_759_im;
    shift_reg_761_re <= shift_reg_760_re;
    shift_reg_761_im <= shift_reg_760_im;
    shift_reg_762_re <= shift_reg_761_re;
    shift_reg_762_im <= shift_reg_761_im;
    shift_reg_763_re <= shift_reg_762_re;
    shift_reg_763_im <= shift_reg_762_im;
    shift_reg_764_re <= shift_reg_763_re;
    shift_reg_764_im <= shift_reg_763_im;
    shift_reg_765_re <= shift_reg_764_re;
    shift_reg_765_im <= shift_reg_764_im;
    shift_reg_766_re <= shift_reg_765_re;
    shift_reg_766_im <= shift_reg_765_im;
    shift_reg_767_re <= shift_reg_766_re;
    shift_reg_767_im <= shift_reg_766_im;
    shift_reg_768_re <= shift_reg_767_re;
    shift_reg_768_im <= shift_reg_767_im;
    shift_reg_769_re <= shift_reg_768_re;
    shift_reg_769_im <= shift_reg_768_im;
    shift_reg_770_re <= shift_reg_769_re;
    shift_reg_770_im <= shift_reg_769_im;
    shift_reg_771_re <= shift_reg_770_re;
    shift_reg_771_im <= shift_reg_770_im;
    shift_reg_772_re <= shift_reg_771_re;
    shift_reg_772_im <= shift_reg_771_im;
    shift_reg_773_re <= shift_reg_772_re;
    shift_reg_773_im <= shift_reg_772_im;
    shift_reg_774_re <= shift_reg_773_re;
    shift_reg_774_im <= shift_reg_773_im;
    shift_reg_775_re <= shift_reg_774_re;
    shift_reg_775_im <= shift_reg_774_im;
    shift_reg_776_re <= shift_reg_775_re;
    shift_reg_776_im <= shift_reg_775_im;
    shift_reg_777_re <= shift_reg_776_re;
    shift_reg_777_im <= shift_reg_776_im;
    shift_reg_778_re <= shift_reg_777_re;
    shift_reg_778_im <= shift_reg_777_im;
    shift_reg_779_re <= shift_reg_778_re;
    shift_reg_779_im <= shift_reg_778_im;
    shift_reg_780_re <= shift_reg_779_re;
    shift_reg_780_im <= shift_reg_779_im;
    shift_reg_781_re <= shift_reg_780_re;
    shift_reg_781_im <= shift_reg_780_im;
    shift_reg_782_re <= shift_reg_781_re;
    shift_reg_782_im <= shift_reg_781_im;
    shift_reg_783_re <= shift_reg_782_re;
    shift_reg_783_im <= shift_reg_782_im;
    shift_reg_784_re <= shift_reg_783_re;
    shift_reg_784_im <= shift_reg_783_im;
    shift_reg_785_re <= shift_reg_784_re;
    shift_reg_785_im <= shift_reg_784_im;
    shift_reg_786_re <= shift_reg_785_re;
    shift_reg_786_im <= shift_reg_785_im;
    shift_reg_787_re <= shift_reg_786_re;
    shift_reg_787_im <= shift_reg_786_im;
    shift_reg_788_re <= shift_reg_787_re;
    shift_reg_788_im <= shift_reg_787_im;
    shift_reg_789_re <= shift_reg_788_re;
    shift_reg_789_im <= shift_reg_788_im;
    shift_reg_790_re <= shift_reg_789_re;
    shift_reg_790_im <= shift_reg_789_im;
    shift_reg_791_re <= shift_reg_790_re;
    shift_reg_791_im <= shift_reg_790_im;
    shift_reg_792_re <= shift_reg_791_re;
    shift_reg_792_im <= shift_reg_791_im;
    shift_reg_793_re <= shift_reg_792_re;
    shift_reg_793_im <= shift_reg_792_im;
    shift_reg_794_re <= shift_reg_793_re;
    shift_reg_794_im <= shift_reg_793_im;
    shift_reg_795_re <= shift_reg_794_re;
    shift_reg_795_im <= shift_reg_794_im;
    shift_reg_796_re <= shift_reg_795_re;
    shift_reg_796_im <= shift_reg_795_im;
    shift_reg_797_re <= shift_reg_796_re;
    shift_reg_797_im <= shift_reg_796_im;
    shift_reg_798_re <= shift_reg_797_re;
    shift_reg_798_im <= shift_reg_797_im;
    shift_reg_799_re <= shift_reg_798_re;
    shift_reg_799_im <= shift_reg_798_im;
    shift_reg_800_re <= shift_reg_799_re;
    shift_reg_800_im <= shift_reg_799_im;
    shift_reg_801_re <= shift_reg_800_re;
    shift_reg_801_im <= shift_reg_800_im;
    shift_reg_802_re <= shift_reg_801_re;
    shift_reg_802_im <= shift_reg_801_im;
    shift_reg_803_re <= shift_reg_802_re;
    shift_reg_803_im <= shift_reg_802_im;
    shift_reg_804_re <= shift_reg_803_re;
    shift_reg_804_im <= shift_reg_803_im;
    shift_reg_805_re <= shift_reg_804_re;
    shift_reg_805_im <= shift_reg_804_im;
    shift_reg_806_re <= shift_reg_805_re;
    shift_reg_806_im <= shift_reg_805_im;
    shift_reg_807_re <= shift_reg_806_re;
    shift_reg_807_im <= shift_reg_806_im;
    shift_reg_808_re <= shift_reg_807_re;
    shift_reg_808_im <= shift_reg_807_im;
    shift_reg_809_re <= shift_reg_808_re;
    shift_reg_809_im <= shift_reg_808_im;
    shift_reg_810_re <= shift_reg_809_re;
    shift_reg_810_im <= shift_reg_809_im;
    shift_reg_811_re <= shift_reg_810_re;
    shift_reg_811_im <= shift_reg_810_im;
    shift_reg_812_re <= shift_reg_811_re;
    shift_reg_812_im <= shift_reg_811_im;
    shift_reg_813_re <= shift_reg_812_re;
    shift_reg_813_im <= shift_reg_812_im;
    shift_reg_814_re <= shift_reg_813_re;
    shift_reg_814_im <= shift_reg_813_im;
    shift_reg_815_re <= shift_reg_814_re;
    shift_reg_815_im <= shift_reg_814_im;
    shift_reg_816_re <= shift_reg_815_re;
    shift_reg_816_im <= shift_reg_815_im;
    shift_reg_817_re <= shift_reg_816_re;
    shift_reg_817_im <= shift_reg_816_im;
    shift_reg_818_re <= shift_reg_817_re;
    shift_reg_818_im <= shift_reg_817_im;
    shift_reg_819_re <= shift_reg_818_re;
    shift_reg_819_im <= shift_reg_818_im;
    shift_reg_820_re <= shift_reg_819_re;
    shift_reg_820_im <= shift_reg_819_im;
    shift_reg_821_re <= shift_reg_820_re;
    shift_reg_821_im <= shift_reg_820_im;
    shift_reg_822_re <= shift_reg_821_re;
    shift_reg_822_im <= shift_reg_821_im;
    shift_reg_823_re <= shift_reg_822_re;
    shift_reg_823_im <= shift_reg_822_im;
    shift_reg_824_re <= shift_reg_823_re;
    shift_reg_824_im <= shift_reg_823_im;
    shift_reg_825_re <= shift_reg_824_re;
    shift_reg_825_im <= shift_reg_824_im;
    shift_reg_826_re <= shift_reg_825_re;
    shift_reg_826_im <= shift_reg_825_im;
    shift_reg_827_re <= shift_reg_826_re;
    shift_reg_827_im <= shift_reg_826_im;
    shift_reg_828_re <= shift_reg_827_re;
    shift_reg_828_im <= shift_reg_827_im;
    shift_reg_829_re <= shift_reg_828_re;
    shift_reg_829_im <= shift_reg_828_im;
    shift_reg_830_re <= shift_reg_829_re;
    shift_reg_830_im <= shift_reg_829_im;
    shift_reg_831_re <= shift_reg_830_re;
    shift_reg_831_im <= shift_reg_830_im;
    shift_reg_832_re <= shift_reg_831_re;
    shift_reg_832_im <= shift_reg_831_im;
    shift_reg_833_re <= shift_reg_832_re;
    shift_reg_833_im <= shift_reg_832_im;
    shift_reg_834_re <= shift_reg_833_re;
    shift_reg_834_im <= shift_reg_833_im;
    shift_reg_835_re <= shift_reg_834_re;
    shift_reg_835_im <= shift_reg_834_im;
    shift_reg_836_re <= shift_reg_835_re;
    shift_reg_836_im <= shift_reg_835_im;
    shift_reg_837_re <= shift_reg_836_re;
    shift_reg_837_im <= shift_reg_836_im;
    shift_reg_838_re <= shift_reg_837_re;
    shift_reg_838_im <= shift_reg_837_im;
    shift_reg_839_re <= shift_reg_838_re;
    shift_reg_839_im <= shift_reg_838_im;
    shift_reg_840_re <= shift_reg_839_re;
    shift_reg_840_im <= shift_reg_839_im;
    shift_reg_841_re <= shift_reg_840_re;
    shift_reg_841_im <= shift_reg_840_im;
    shift_reg_842_re <= shift_reg_841_re;
    shift_reg_842_im <= shift_reg_841_im;
    shift_reg_843_re <= shift_reg_842_re;
    shift_reg_843_im <= shift_reg_842_im;
    shift_reg_844_re <= shift_reg_843_re;
    shift_reg_844_im <= shift_reg_843_im;
    shift_reg_845_re <= shift_reg_844_re;
    shift_reg_845_im <= shift_reg_844_im;
    shift_reg_846_re <= shift_reg_845_re;
    shift_reg_846_im <= shift_reg_845_im;
    shift_reg_847_re <= shift_reg_846_re;
    shift_reg_847_im <= shift_reg_846_im;
    shift_reg_848_re <= shift_reg_847_re;
    shift_reg_848_im <= shift_reg_847_im;
    shift_reg_849_re <= shift_reg_848_re;
    shift_reg_849_im <= shift_reg_848_im;
    shift_reg_850_re <= shift_reg_849_re;
    shift_reg_850_im <= shift_reg_849_im;
    shift_reg_851_re <= shift_reg_850_re;
    shift_reg_851_im <= shift_reg_850_im;
    shift_reg_852_re <= shift_reg_851_re;
    shift_reg_852_im <= shift_reg_851_im;
    shift_reg_853_re <= shift_reg_852_re;
    shift_reg_853_im <= shift_reg_852_im;
    shift_reg_854_re <= shift_reg_853_re;
    shift_reg_854_im <= shift_reg_853_im;
    shift_reg_855_re <= shift_reg_854_re;
    shift_reg_855_im <= shift_reg_854_im;
    shift_reg_856_re <= shift_reg_855_re;
    shift_reg_856_im <= shift_reg_855_im;
    shift_reg_857_re <= shift_reg_856_re;
    shift_reg_857_im <= shift_reg_856_im;
    shift_reg_858_re <= shift_reg_857_re;
    shift_reg_858_im <= shift_reg_857_im;
    shift_reg_859_re <= shift_reg_858_re;
    shift_reg_859_im <= shift_reg_858_im;
    shift_reg_860_re <= shift_reg_859_re;
    shift_reg_860_im <= shift_reg_859_im;
    shift_reg_861_re <= shift_reg_860_re;
    shift_reg_861_im <= shift_reg_860_im;
    shift_reg_862_re <= shift_reg_861_re;
    shift_reg_862_im <= shift_reg_861_im;
    shift_reg_863_re <= shift_reg_862_re;
    shift_reg_863_im <= shift_reg_862_im;
    shift_reg_864_re <= shift_reg_863_re;
    shift_reg_864_im <= shift_reg_863_im;
    shift_reg_865_re <= shift_reg_864_re;
    shift_reg_865_im <= shift_reg_864_im;
    shift_reg_866_re <= shift_reg_865_re;
    shift_reg_866_im <= shift_reg_865_im;
    shift_reg_867_re <= shift_reg_866_re;
    shift_reg_867_im <= shift_reg_866_im;
    shift_reg_868_re <= shift_reg_867_re;
    shift_reg_868_im <= shift_reg_867_im;
    shift_reg_869_re <= shift_reg_868_re;
    shift_reg_869_im <= shift_reg_868_im;
    shift_reg_870_re <= shift_reg_869_re;
    shift_reg_870_im <= shift_reg_869_im;
    shift_reg_871_re <= shift_reg_870_re;
    shift_reg_871_im <= shift_reg_870_im;
    shift_reg_872_re <= shift_reg_871_re;
    shift_reg_872_im <= shift_reg_871_im;
    shift_reg_873_re <= shift_reg_872_re;
    shift_reg_873_im <= shift_reg_872_im;
    shift_reg_874_re <= shift_reg_873_re;
    shift_reg_874_im <= shift_reg_873_im;
    shift_reg_875_re <= shift_reg_874_re;
    shift_reg_875_im <= shift_reg_874_im;
    shift_reg_876_re <= shift_reg_875_re;
    shift_reg_876_im <= shift_reg_875_im;
    shift_reg_877_re <= shift_reg_876_re;
    shift_reg_877_im <= shift_reg_876_im;
    shift_reg_878_re <= shift_reg_877_re;
    shift_reg_878_im <= shift_reg_877_im;
    shift_reg_879_re <= shift_reg_878_re;
    shift_reg_879_im <= shift_reg_878_im;
    shift_reg_880_re <= shift_reg_879_re;
    shift_reg_880_im <= shift_reg_879_im;
    shift_reg_881_re <= shift_reg_880_re;
    shift_reg_881_im <= shift_reg_880_im;
    shift_reg_882_re <= shift_reg_881_re;
    shift_reg_882_im <= shift_reg_881_im;
    shift_reg_883_re <= shift_reg_882_re;
    shift_reg_883_im <= shift_reg_882_im;
    shift_reg_884_re <= shift_reg_883_re;
    shift_reg_884_im <= shift_reg_883_im;
    shift_reg_885_re <= shift_reg_884_re;
    shift_reg_885_im <= shift_reg_884_im;
    shift_reg_886_re <= shift_reg_885_re;
    shift_reg_886_im <= shift_reg_885_im;
    shift_reg_887_re <= shift_reg_886_re;
    shift_reg_887_im <= shift_reg_886_im;
    shift_reg_888_re <= shift_reg_887_re;
    shift_reg_888_im <= shift_reg_887_im;
    shift_reg_889_re <= shift_reg_888_re;
    shift_reg_889_im <= shift_reg_888_im;
    shift_reg_890_re <= shift_reg_889_re;
    shift_reg_890_im <= shift_reg_889_im;
    shift_reg_891_re <= shift_reg_890_re;
    shift_reg_891_im <= shift_reg_890_im;
    shift_reg_892_re <= shift_reg_891_re;
    shift_reg_892_im <= shift_reg_891_im;
    shift_reg_893_re <= shift_reg_892_re;
    shift_reg_893_im <= shift_reg_892_im;
    shift_reg_894_re <= shift_reg_893_re;
    shift_reg_894_im <= shift_reg_893_im;
    shift_reg_895_re <= shift_reg_894_re;
    shift_reg_895_im <= shift_reg_894_im;
    shift_reg_896_re <= shift_reg_895_re;
    shift_reg_896_im <= shift_reg_895_im;
    shift_reg_897_re <= shift_reg_896_re;
    shift_reg_897_im <= shift_reg_896_im;
    shift_reg_898_re <= shift_reg_897_re;
    shift_reg_898_im <= shift_reg_897_im;
    shift_reg_899_re <= shift_reg_898_re;
    shift_reg_899_im <= shift_reg_898_im;
    shift_reg_900_re <= shift_reg_899_re;
    shift_reg_900_im <= shift_reg_899_im;
    shift_reg_901_re <= shift_reg_900_re;
    shift_reg_901_im <= shift_reg_900_im;
    shift_reg_902_re <= shift_reg_901_re;
    shift_reg_902_im <= shift_reg_901_im;
    shift_reg_903_re <= shift_reg_902_re;
    shift_reg_903_im <= shift_reg_902_im;
    shift_reg_904_re <= shift_reg_903_re;
    shift_reg_904_im <= shift_reg_903_im;
    shift_reg_905_re <= shift_reg_904_re;
    shift_reg_905_im <= shift_reg_904_im;
    shift_reg_906_re <= shift_reg_905_re;
    shift_reg_906_im <= shift_reg_905_im;
    shift_reg_907_re <= shift_reg_906_re;
    shift_reg_907_im <= shift_reg_906_im;
    shift_reg_908_re <= shift_reg_907_re;
    shift_reg_908_im <= shift_reg_907_im;
    shift_reg_909_re <= shift_reg_908_re;
    shift_reg_909_im <= shift_reg_908_im;
    shift_reg_910_re <= shift_reg_909_re;
    shift_reg_910_im <= shift_reg_909_im;
    shift_reg_911_re <= shift_reg_910_re;
    shift_reg_911_im <= shift_reg_910_im;
    shift_reg_912_re <= shift_reg_911_re;
    shift_reg_912_im <= shift_reg_911_im;
    shift_reg_913_re <= shift_reg_912_re;
    shift_reg_913_im <= shift_reg_912_im;
    shift_reg_914_re <= shift_reg_913_re;
    shift_reg_914_im <= shift_reg_913_im;
    shift_reg_915_re <= shift_reg_914_re;
    shift_reg_915_im <= shift_reg_914_im;
    shift_reg_916_re <= shift_reg_915_re;
    shift_reg_916_im <= shift_reg_915_im;
    shift_reg_917_re <= shift_reg_916_re;
    shift_reg_917_im <= shift_reg_916_im;
    shift_reg_918_re <= shift_reg_917_re;
    shift_reg_918_im <= shift_reg_917_im;
    shift_reg_919_re <= shift_reg_918_re;
    shift_reg_919_im <= shift_reg_918_im;
    shift_reg_920_re <= shift_reg_919_re;
    shift_reg_920_im <= shift_reg_919_im;
    shift_reg_921_re <= shift_reg_920_re;
    shift_reg_921_im <= shift_reg_920_im;
    shift_reg_922_re <= shift_reg_921_re;
    shift_reg_922_im <= shift_reg_921_im;
    shift_reg_923_re <= shift_reg_922_re;
    shift_reg_923_im <= shift_reg_922_im;
    shift_reg_924_re <= shift_reg_923_re;
    shift_reg_924_im <= shift_reg_923_im;
    shift_reg_925_re <= shift_reg_924_re;
    shift_reg_925_im <= shift_reg_924_im;
    shift_reg_926_re <= shift_reg_925_re;
    shift_reg_926_im <= shift_reg_925_im;
    shift_reg_927_re <= shift_reg_926_re;
    shift_reg_927_im <= shift_reg_926_im;
    shift_reg_928_re <= shift_reg_927_re;
    shift_reg_928_im <= shift_reg_927_im;
    shift_reg_929_re <= shift_reg_928_re;
    shift_reg_929_im <= shift_reg_928_im;
    shift_reg_930_re <= shift_reg_929_re;
    shift_reg_930_im <= shift_reg_929_im;
    shift_reg_931_re <= shift_reg_930_re;
    shift_reg_931_im <= shift_reg_930_im;
    shift_reg_932_re <= shift_reg_931_re;
    shift_reg_932_im <= shift_reg_931_im;
    shift_reg_933_re <= shift_reg_932_re;
    shift_reg_933_im <= shift_reg_932_im;
    shift_reg_934_re <= shift_reg_933_re;
    shift_reg_934_im <= shift_reg_933_im;
    shift_reg_935_re <= shift_reg_934_re;
    shift_reg_935_im <= shift_reg_934_im;
    shift_reg_936_re <= shift_reg_935_re;
    shift_reg_936_im <= shift_reg_935_im;
    shift_reg_937_re <= shift_reg_936_re;
    shift_reg_937_im <= shift_reg_936_im;
    shift_reg_938_re <= shift_reg_937_re;
    shift_reg_938_im <= shift_reg_937_im;
    shift_reg_939_re <= shift_reg_938_re;
    shift_reg_939_im <= shift_reg_938_im;
    shift_reg_940_re <= shift_reg_939_re;
    shift_reg_940_im <= shift_reg_939_im;
    shift_reg_941_re <= shift_reg_940_re;
    shift_reg_941_im <= shift_reg_940_im;
    shift_reg_942_re <= shift_reg_941_re;
    shift_reg_942_im <= shift_reg_941_im;
    shift_reg_943_re <= shift_reg_942_re;
    shift_reg_943_im <= shift_reg_942_im;
    shift_reg_944_re <= shift_reg_943_re;
    shift_reg_944_im <= shift_reg_943_im;
    shift_reg_945_re <= shift_reg_944_re;
    shift_reg_945_im <= shift_reg_944_im;
    shift_reg_946_re <= shift_reg_945_re;
    shift_reg_946_im <= shift_reg_945_im;
    shift_reg_947_re <= shift_reg_946_re;
    shift_reg_947_im <= shift_reg_946_im;
    shift_reg_948_re <= shift_reg_947_re;
    shift_reg_948_im <= shift_reg_947_im;
    shift_reg_949_re <= shift_reg_948_re;
    shift_reg_949_im <= shift_reg_948_im;
    shift_reg_950_re <= shift_reg_949_re;
    shift_reg_950_im <= shift_reg_949_im;
    shift_reg_951_re <= shift_reg_950_re;
    shift_reg_951_im <= shift_reg_950_im;
    shift_reg_952_re <= shift_reg_951_re;
    shift_reg_952_im <= shift_reg_951_im;
    shift_reg_953_re <= shift_reg_952_re;
    shift_reg_953_im <= shift_reg_952_im;
    shift_reg_954_re <= shift_reg_953_re;
    shift_reg_954_im <= shift_reg_953_im;
    shift_reg_955_re <= shift_reg_954_re;
    shift_reg_955_im <= shift_reg_954_im;
    shift_reg_956_re <= shift_reg_955_re;
    shift_reg_956_im <= shift_reg_955_im;
    shift_reg_957_re <= shift_reg_956_re;
    shift_reg_957_im <= shift_reg_956_im;
    shift_reg_958_re <= shift_reg_957_re;
    shift_reg_958_im <= shift_reg_957_im;
    shift_reg_959_re <= shift_reg_958_re;
    shift_reg_959_im <= shift_reg_958_im;
    shift_reg_960_re <= shift_reg_959_re;
    shift_reg_960_im <= shift_reg_959_im;
    shift_reg_961_re <= shift_reg_960_re;
    shift_reg_961_im <= shift_reg_960_im;
    shift_reg_962_re <= shift_reg_961_re;
    shift_reg_962_im <= shift_reg_961_im;
    shift_reg_963_re <= shift_reg_962_re;
    shift_reg_963_im <= shift_reg_962_im;
    shift_reg_964_re <= shift_reg_963_re;
    shift_reg_964_im <= shift_reg_963_im;
    shift_reg_965_re <= shift_reg_964_re;
    shift_reg_965_im <= shift_reg_964_im;
    shift_reg_966_re <= shift_reg_965_re;
    shift_reg_966_im <= shift_reg_965_im;
    shift_reg_967_re <= shift_reg_966_re;
    shift_reg_967_im <= shift_reg_966_im;
    shift_reg_968_re <= shift_reg_967_re;
    shift_reg_968_im <= shift_reg_967_im;
    shift_reg_969_re <= shift_reg_968_re;
    shift_reg_969_im <= shift_reg_968_im;
    shift_reg_970_re <= shift_reg_969_re;
    shift_reg_970_im <= shift_reg_969_im;
    shift_reg_971_re <= shift_reg_970_re;
    shift_reg_971_im <= shift_reg_970_im;
    shift_reg_972_re <= shift_reg_971_re;
    shift_reg_972_im <= shift_reg_971_im;
    shift_reg_973_re <= shift_reg_972_re;
    shift_reg_973_im <= shift_reg_972_im;
    shift_reg_974_re <= shift_reg_973_re;
    shift_reg_974_im <= shift_reg_973_im;
    shift_reg_975_re <= shift_reg_974_re;
    shift_reg_975_im <= shift_reg_974_im;
    shift_reg_976_re <= shift_reg_975_re;
    shift_reg_976_im <= shift_reg_975_im;
    shift_reg_977_re <= shift_reg_976_re;
    shift_reg_977_im <= shift_reg_976_im;
    shift_reg_978_re <= shift_reg_977_re;
    shift_reg_978_im <= shift_reg_977_im;
    shift_reg_979_re <= shift_reg_978_re;
    shift_reg_979_im <= shift_reg_978_im;
    shift_reg_980_re <= shift_reg_979_re;
    shift_reg_980_im <= shift_reg_979_im;
    shift_reg_981_re <= shift_reg_980_re;
    shift_reg_981_im <= shift_reg_980_im;
    shift_reg_982_re <= shift_reg_981_re;
    shift_reg_982_im <= shift_reg_981_im;
    shift_reg_983_re <= shift_reg_982_re;
    shift_reg_983_im <= shift_reg_982_im;
    shift_reg_984_re <= shift_reg_983_re;
    shift_reg_984_im <= shift_reg_983_im;
    shift_reg_985_re <= shift_reg_984_re;
    shift_reg_985_im <= shift_reg_984_im;
    shift_reg_986_re <= shift_reg_985_re;
    shift_reg_986_im <= shift_reg_985_im;
    shift_reg_987_re <= shift_reg_986_re;
    shift_reg_987_im <= shift_reg_986_im;
    shift_reg_988_re <= shift_reg_987_re;
    shift_reg_988_im <= shift_reg_987_im;
    shift_reg_989_re <= shift_reg_988_re;
    shift_reg_989_im <= shift_reg_988_im;
    shift_reg_990_re <= shift_reg_989_re;
    shift_reg_990_im <= shift_reg_989_im;
    shift_reg_991_re <= shift_reg_990_re;
    shift_reg_991_im <= shift_reg_990_im;
    shift_reg_992_re <= shift_reg_991_re;
    shift_reg_992_im <= shift_reg_991_im;
    shift_reg_993_re <= shift_reg_992_re;
    shift_reg_993_im <= shift_reg_992_im;
    shift_reg_994_re <= shift_reg_993_re;
    shift_reg_994_im <= shift_reg_993_im;
    shift_reg_995_re <= shift_reg_994_re;
    shift_reg_995_im <= shift_reg_994_im;
    shift_reg_996_re <= shift_reg_995_re;
    shift_reg_996_im <= shift_reg_995_im;
    shift_reg_997_re <= shift_reg_996_re;
    shift_reg_997_im <= shift_reg_996_im;
    shift_reg_998_re <= shift_reg_997_re;
    shift_reg_998_im <= shift_reg_997_im;
    shift_reg_999_re <= shift_reg_998_re;
    shift_reg_999_im <= shift_reg_998_im;
    shift_reg_1000_re <= shift_reg_999_re;
    shift_reg_1000_im <= shift_reg_999_im;
    shift_reg_1001_re <= shift_reg_1000_re;
    shift_reg_1001_im <= shift_reg_1000_im;
    shift_reg_1002_re <= shift_reg_1001_re;
    shift_reg_1002_im <= shift_reg_1001_im;
    shift_reg_1003_re <= shift_reg_1002_re;
    shift_reg_1003_im <= shift_reg_1002_im;
    shift_reg_1004_re <= shift_reg_1003_re;
    shift_reg_1004_im <= shift_reg_1003_im;
    shift_reg_1005_re <= shift_reg_1004_re;
    shift_reg_1005_im <= shift_reg_1004_im;
    shift_reg_1006_re <= shift_reg_1005_re;
    shift_reg_1006_im <= shift_reg_1005_im;
    shift_reg_1007_re <= shift_reg_1006_re;
    shift_reg_1007_im <= shift_reg_1006_im;
    shift_reg_1008_re <= shift_reg_1007_re;
    shift_reg_1008_im <= shift_reg_1007_im;
    shift_reg_1009_re <= shift_reg_1008_re;
    shift_reg_1009_im <= shift_reg_1008_im;
    shift_reg_1010_re <= shift_reg_1009_re;
    shift_reg_1010_im <= shift_reg_1009_im;
    shift_reg_1011_re <= shift_reg_1010_re;
    shift_reg_1011_im <= shift_reg_1010_im;
    shift_reg_1012_re <= shift_reg_1011_re;
    shift_reg_1012_im <= shift_reg_1011_im;
    shift_reg_1013_re <= shift_reg_1012_re;
    shift_reg_1013_im <= shift_reg_1012_im;
    shift_reg_1014_re <= shift_reg_1013_re;
    shift_reg_1014_im <= shift_reg_1013_im;
    shift_reg_1015_re <= shift_reg_1014_re;
    shift_reg_1015_im <= shift_reg_1014_im;
    shift_reg_1016_re <= shift_reg_1015_re;
    shift_reg_1016_im <= shift_reg_1015_im;
    shift_reg_1017_re <= shift_reg_1016_re;
    shift_reg_1017_im <= shift_reg_1016_im;
    shift_reg_1018_re <= shift_reg_1017_re;
    shift_reg_1018_im <= shift_reg_1017_im;
    shift_reg_1019_re <= shift_reg_1018_re;
    shift_reg_1019_im <= shift_reg_1018_im;
    shift_reg_1020_re <= shift_reg_1019_re;
    shift_reg_1020_im <= shift_reg_1019_im;
    shift_reg_1021_re <= shift_reg_1020_re;
    shift_reg_1021_im <= shift_reg_1020_im;
    shift_reg_1022_re <= shift_reg_1021_re;
    shift_reg_1022_im <= shift_reg_1021_im;
    shift_reg_1023_re <= shift_reg_1022_re;
    shift_reg_1023_im <= shift_reg_1022_im;
  end


endmodule
